även i vår värld finns floder och träd och lejon och elefanter .
står upp , går till ett hörn , den skälver ,
Historien jag har berättat för er är stökig och oavslutad .
central Intelligence Agency .
Låt oss leva med varandra och ta ett andetag i taget .
det är en gentleman på första raden som faktiskt gör en exakt imitation av hur hon såg ut .
vi vinner mark och snart kommer vi att övervinna krisen .
hos de här barnen ville jag föra tanken till något som existerar inombords som ingen kan ta bort , så jag utarbetade en kursplan som dels är statsvetenskap , dels fotbollsturnering , i en konstfestival .
det beklagliga är att våra städer , som New Delhi och Mumbai , inte har tillgång till vatten dygnet runt .
ni kan om ni vill jämföra detta med , å ena sidan en hjärtinfarkt där man har död vävnad i hjärtat , kontra arytmi , där ett organ helt enkelt inte fungerar på grund av kommunikationsproblem inuti det .
om du är ogift , sjunker siffran till tre .
så detta är vad vi kallar en oktaeder .
innan jag går vidare vill jag förtydliga min egen roll i detta .
vi tog en annan grupp , en stor grupp amerikaner , och ställde en fråga i okunnighetens slöja .
men , jag vet själv också , jag känner den här virtuella esprit de corps , om ni så vill , med dem allihop .
vad pågår i den här bebisens huvud ?
kaffe både orsakar och motverkar cancer .
den uppenbara frågan är , behöver verkligen ett TEDTalk 2300 ord ?
( Applåder ) ca : under tiden , med hjälp av internet och den här tekniken , är du här , tillbaka i Nordamerika , inte riktigt USA , men Kanada , på det här sättet .
verkligen inte . Låt oss se till att de närmsta 100 åren blir det bästa av århundraden .
nummer 5 : Osäkerhetsmomentet .
jag skrev den här efter en väns begravning men inte så mycket om vännen som om något griftetalaren pratade om som alla griftetalare brukar göra , vilket är hur glad den avlidne skulle varit om hen tittade ner och såg oss alla samlade .
Doktor King trodde på att de fanns två typer av lagar i denna värld , de som skapas av en högre makt och de som skapas av människor .
du ska till sydamerika , inte sant ? &quot;
( Skratt ) Om jag går för långt åt andra hållet och gör det väldigt abstrakt vet ingen vad det är de ser .
det här kanske ligger på gränsen till science fiction , men om även en liten del av det här scenariot blir sanning kommer vår ekologi och till och med vår art inte att klara sig länge oskadda ifrån det .
så allt jag stoppade i min kropp ansåg jag vara medicin .
ett av testen vi använde för kreativitet var alternativa användningsområden .
jag arbetar med morgondagens forskare och ledare , och de förtjänar att få reda på vad vetenskapen säger så att de kan hjälpa till att forma en framtid för alla .
Beteendeekonomen Georg Lowenstein bad studenter på sitt universitet föreställa sig att få en passionerad kyss från en berömd person , vilken som helst .
den var beviset på att jag inte hade räckt till , att jag var gammal och inte fantastisk och inte perfekt och inte passade in i den förutbestämda mallen .
jag vet inget annat om honom , utom att han en gång räddade mitt liv genom att riskera sitt eget .
vi behöver kunna säga någonting , för vet ni vilka fler som sitter vid bordet ?
han lyckades få till ett möte med fader Samaan , och överraskande nog älskade han idén .
du ser att de som väntar till sista minuten har så fullt upp med annat att de inte har några nya idéer .
men det provades aldrig .
kära föräldrar , om ni skäms för mens , så kommer era döttrar göra det också .
svar : det tog dem , i genomsnitt , tre och en halv minut längre tid .
och det är endast när vi hedrar dem och uppmärksammar dem och ger dem status som världen verkligen kommer att förändras .
jag kom bara på besök och sade , &quot; Det ser bra ut , bra jobbat &quot; , Det var allt . ni kan se vad klockan är i alla fem kommuner av New York där bak . så det här är utrymmet för handledningstimmarna .
( Skratt ) och en man kom att ge berättelser om sin far genom en plattform som heter Twitter för att kommunicera den skit hans far kom att uttrycka .
det var en ordentlig utmaning , och det var faktiskt exempel från biologi som bidrog oss med många av ledtrådarna .
varför vi väljer de semestrar vi väljer är ett problem vi möter med ett val mellan de två själven .
och farmor , var fanns du när de marscherade med våra japansk @-@ amerikanska grannar till interneringslägren ?
så låg inkomst här och hög inkomst här .
på andra områden snöar det eller så ökar ismassan igen på vintern .
och om människor flyttar till urbana , okända , betongmiljöer så kan de också bli hjälpta i förväg av socialt stöd som redan väntar genom SMS @-@ kunskap .
trots det , 70 år senare , har cirkeln slutits .
och i denna stund är vi perfekta , vi är hela och vi är vackra .
Bryr vi oss om människorna , vår familj , hälsa , eller är det prestation , framgång , sådant ?
Sömnkvaliteten som du får som nattskiftsarbetare är normalt sett mycket dålig , återigen i femtimmarsregionen .
det betyder inte att vi nödvändigtvis kommer till samma slutsats .
han hade en mycket generös returpolicy , detaljerade köpvillkor , och kort leveranstid .
och nu ska vi tända på det .
en dollar , tio dollar eller 100 dollar per dag .
så snart den tilliten var uppbyggd ville alla vara med på vårt maraton för att visa världen Libanons sanna färger och det Libanesiska folket och deras önskan att leva i fred och harmoni .
små finjusteringar kan leda till stora förändringar .
så jag hoppas ni gillar det .
det använder inte optik som ett vanligt mikroskop för att göra små objekt större . Istället använder den en videokamera och bildbehandling för att avslöja de minsta rörelserna och färgförändringarna hos saker och människor förändringar som är omöjliga för oss att se med blotta ögat ,
nu ser vi en stark ökning av nya konflikter och de gamla konflikterna är kvar : Afganistan , Somalia , demokratiska republiken Kongo .
jag var så hänförd av resultatet att jag ville plantera dessa skogar på samma sätt som vi tillverkar bilar , skriver programvara , eller driver vanliga verksamheter , så jag grundade ett företag , en end @-@ To @-@ end tjänst , för att skapa dessa inhemska naturskogar .
med den här inställningen . den andra aspekten av min livsfilosofi är att jag omger mig med människor som jag vill vara med , människor av god kvalitet .
vad alla dessa människor har gemensamt är att de är kättare .
Lunginflammation tog tre barn av tio .
ta till exempel Airbnbs massiva succé som alla känner till .
i intervjun pratar hon med sin dotter Lesley om att som ung man gå med i ett gäng , och senare i livet bli den kvinna hon alltid var ämnad att bli .
för 150 år sedan beskrev anatomer väldigt , väldigt noggrant -- här har ni en modell av magväggen .
när en fluga rör sig över mittpunkten i kammaren där de två strömmarna av luktämnen möts , måste den ta ett beslut .
och ingen skulle ge sitt livs besparingar till ökända smugglare om det fanns en laglig väg för migration .
Utförandezonen maximerar våra omedelbara resultat , och inlärningszonen vår utveckling och framtida prestation .
och en sak man ser är att på manslinjen går dödligheten neråt , neråt , neråt , neråt , neråt .
det var frihet under ansvar .
innan vaccinerna fanns dödade många av infektionssjukdomarna miljontals människor per år .
och det är mycket mer på gång .
hon ville skapa ett bättre liv för sina barn och sin familj .
om du verkligen bryr dig om att starta en rörelse , ha modet att följa och att visa andra hur man följer .
de är också silikon .
jag är här för att berätta för er om framgång i Afrika .
men finns det tänkbara händelser som kan vara ännu värre , som kan släcka ut allt liv ?
hur många av er använder skrivbordsfältet ?
Undersökningsrummet kändes som ett skämt .
PM : det tror jag inte . NA : men det hjälper att berätta att några människor är agenter för förändring i samhället .
som den där spindeln som bor bakom din soffa ?
men det är fortfarande lite komplicerat och lite svårt .
mitt företag har mjukvara som gör detta redan idag .
tack så mycket , Chris .
jag undrade om vi kunde använda all data och all vår expertkunskap när vi utvecklar nätverk för att kvantifiera hur detta kan ske .
men okej är aldrig okej .
för att nummer ett , svaret spelar roll .
varje land i världen har tidningar . den har ett bisarrt på pågående filosofisk projekt ,
så människor går omkring med virus som inte märks .
dessa barn växer upp utan familjeförebilder eller en bild av goda föräldrar , så de kan ha svårt att själva vara föräldrar åt sina egna barn .
detta är en plats av stor historisk betydelse .
och om du drar på den här sidan av repet , försvinner repet från den andra sidan .
vi ska inte oroa oss för vad våra maskiner kan göra idag .
vi åkte tillbaka för den sista visningen av gården , och han visade mig de vilda pepparplantorna och växterna som han såg till fanns där för sältan .
Vår framtid är många @-@ till @-@ många .
Nyfikenhet och förundran , för den driver oss att utforska , för vi är omgivna av saker som vi inte kan se .
det finns ingen som inte har gjort det så här långt .
det är de blå staplarna .
det var för fem år sen som jag verkligen började bryta ny mark genom att kombinera virtual reality och journalistik .
så häng med mig runt och tillbaka i resonemanget .
och det ledde sedan till Mina stora frågor .
Ammoniaken avdunstar och den återkondenserar på andra sidan .
just nu kan datorer göra det som människor ägnar det mesta av sin tid åt att göra för att få betalt , så det är hög tid att börja tänka på hur vi ska anpassa våra sociala och ekonomiska strukturer för att klara av den nya verkligheten .
trots det är dessa miljöer bra platser för att stoppa den rörliga sanden .
det förändrar hur du hanterar din upplevelse , det förändrar hur du tänker på din förövare , det betyder att om du träder fram , backar du upp någon annan och de backar upp dig .
så livet måste förändras .
så jag sprang ut i vinterkylan och fotograferade varenda person jag kunde få tag på i februari för två år sedan .
lokal jihad blir Global jihad igen om man struntar i det .
hur löser då hjärnan sitt avfallsproblem ?
han fick sin arm amputerad för 10 år sedan .
och vi beslöt att vi på minsta möjliga tid skulle förstå hur det nya viruset betedde sig i våra barn .
( Maskinröst ) 1,8 . vi har många försök igång ute i byarna och i skolorna , och utifrån vad vi lärt oss ute i fält , har vi insett att det är viktigt att använda icke @-@ medicinska termer så att människor kan förstå vad vi undersöker och vad det betyder för dem .
och det verkar vara ett tryggt levnadssätt .
så , på grund av den här explosionen i ljudtillgänglighet särskilt hos döva har detta inte bara påverkat hur musikinstitutioner och dövskolor behandlar ljud - och inte bara som terapimetod - fast som medgestaltare av musik , stämmer detta absolut också . men det har betytt att akustiker verkligen har behövt fundera över vilka slags lokaler de konstruerar .
flera år efter denna händelse tränade han racketbolltränarna .
för jag är kvinna .
men en fantastisk person var han , en underbar filosof .
det är en av de saker jag är mest stolt över i mitt liv .
Publiken : 23
så jag säger till honom , helt klart i mitt huvud : &quot; det är Jill , jag behöver hjälp ! &quot;
när vi letar upp dem och frågar vad det är så säger de oftast något i stil med : &quot; jag är helt enkelt inte någon kreativ person &quot; .
och när hon växte upp , när hon var fyra och ett halvt år gammal , skrev jag in henne i min skola .
en tid efter att den kom ut , väntade Augusten på en flygplats och besökte bokhandeln och tittade på vilka som köpte hans böcker .
jag började med det för 15 år sen .
och sen kom killen på en briljant idé , han sa , &quot; Du driver ju den där organisationen ungdomar utan gränser , eller hur ?
så jag tog reda på vad ekonomin betalade för kriget i Irak samma år .
som många andra lägger jag mycket tid på att klaga över hur svårt det är att få människor att förändras , och vi borde inte tjafsa om det .
för när det gäller sex , är män pressade till att skryta och överdriva , medan kvinnor är pressade till att dölja , förminska och förneka , vilket inte är konstigt när man tänker på att det fortfarande finns nio länder där kvinnor kan avrättas för att de vänsterprasslar .
förra året lyckades vi dock skrapa ihop lite pengar .
( Skratt ) ( Applåder ) När vinden blåser , leds all överskottsenergi från vindkraftverket om till batteriet .
att återta våra berättelser och lyssna på varandras , kan skapa en portal som kan överträffa tiden självt .
som tur är så har vi en ny maskin , magnetencefalografi , som låter oss göra detta .
Uppmärksamhet är valutan .
vi ser ett tydligt behov av att aktivt främja hälsoinsatser , särskilt bland äldre .
jag har funderat och vägt samman hur det är att arbeta under kapitalism .
när han gör så , betyder det inte &quot; ta din Stradivarius och som Jimi Hendrix , slå den mot golvet &quot; .
Kometen är alltså fräsch och ny .
det finns andra som nästan faller ihop när de kommer in , man ser det .
var var den här för 10 år sen ?
folk vill alltid berätta saker om sina fantastiska skor .
ändå spenderar vi överraskande lite tid för att ta hand om det som betyder mest : sättet vårt medvetande fungerar . vilket , återigen , är det avgörande som avgör kvalitén på vad vi upplever .
när vi lär känna någon , lär vi oss hur de fungerar , och sedan lär vi oss vilka ämnen vi kan prata om .
då kan vi börja använda celler .
Flickorna själva såg aldrig bilderna , men de gav dem till oss . det är detta som kritikerna inte känner till , och det är denna forskning jag rekommenderar för de som vill arbeta humanistiskt .
hon skulle antagligen säga att hon inte är så speciell , men hon har ett märkvärdigt inflytande .
och , till skillnad från en massa choklad , kan massor av leenden faktisk göra dig friskare .
det var inte okunnighet .
jag var klar med skolan och skulle arbeta som juridiskt ombud och representera stammar runtom i landet , representera på Capitol Hill , och jag såg direkt varför rasistiskt bildspråk spelar roll .
Imorgon kommer det inte finnas någon ursäkt för att inte göra det rätta .
och jag säger er att detta inte är en fråga om klimatpolitik eller miljöpolitik .
och jag tänkte , jag ger dem ett prov . de kommer att få en nolla . sen ger jag dem materialet . jag kommer tillbaka och testar dem . de får en till nolla . och går tillbaka tillbaka och säger , &quot; ja , vi behöver lärare för vissa saker &quot; .
så fort som vi - och detta var på 50 @-@ talet - och så fort som vi tog bort det jagande , trummslagande folket för att skydda djuren , så började marken att försämras , som ni ser i den här parken vi skapade .
så vi började prata om det här .
detsamma är sant för genomskinliga solceller som är integrerade med fönster , solceller integrerade med gatumöbler , eller solceller integrerade med dessa miljarder apparater som bildar Sakernas Internet .
till vänster har vi Casablanca , till höger har vi Chicago .
om vi äter otillagad mat kan vi inte frigöra energin ordentligt .
kort sagt spelar jag in en sekund av mitt liv varje dag i resten av mitt liv , och sedan i tidsordning sätta ihop alla dessa pyttesmå en @-@ sekundare av mitt liv till en lång video tills jag liksom inte kan spela in längre .
jag svarar , &quot; Var inte oroliga , era föräldrar kan inte heller .
ni känner alla till den här historien .
när män säger det handlar det ofta om något som de inte skulle ha gjort ändå .
man filmar vägskyltar , klockor , dagstidningar .
Låt oss till exempel anta att det första fallet inträffar i Sydasien .
det är inget fel på din hjärna . det är inget fel på ditt förstånd . du har Charles Bonnet @-@ syndrom &quot;
Revolutionen inom dödsvård har börjat .
Istället för att säga att det handlar om att vinna tävlingen , kommer folk inse att framgång mer handlar om att bidra .
och uppfinningsrikedomen , om du nu kan kalla det för det , går djupare än så .
det ligger på 826 Valencia Street i Mission @-@ området i San Francisco , och när jag jobbade där låg högkvarteret för ett bokförlag där , som hette McSweeney &apos; s ; en ideell skrivverkstad som hette 826 Valencia . Längst fram i huset låg en märklig affär .
den använder de senaste molekylärbiologiska rönen , och är en billig , 3D @-@ printad enhet , och datavetenskap för att försöka tackla en av mänsklighetens svåraste utmaningar .
och hon bara : - Haha , något sådant finns inte .
i filmen &quot; Spirited away &quot; råkar de som tar emot guld från No @-@ Face ut för otur .
hon väntade otåligt på att flytta hemifrån. för att bevisa för dem att hon är vuxen , och för att bevisa för sina nya vänner att hon är en av dem .
Barnäktenskapen kommer kanske inte att bli färre .
han är någon som flydde från allt detta dåliga &quot; .
det är ett ställe vi går till för att komma bort från stressen i arbetslivet och ibland i familjelivet .
på franska till exempel skulle man säga &quot; tu &quot; när man pratar med sin kompis i skolan men &quot; vous &quot; när man pratar med sin lärare .
det ni alla gör just nu med er bröstkorg , och sluta inte göra det , är att andas . man använder interkostalmusklerna , musklerna mellan revbenen
och deras kunder och miljön .
vi följer dem som leder , inte för deras skull , men för oss vår egen skull .
Arkitekturens välbeprövade och genomtänkta formler och termer fungerar inte här .
som resultat , tycker jag att vi stackars förtryckta kvinnor faktiskt har några nyttiga , surt förvärvade lärdomar att lära ut , lärdomar som kan visa sig användbara för den som vill blomstra i den moderna världen .
IndiGenomics handlar om vetenskap för folket och av folket .
jag blev kallad en idiot , en förrädare , ett plågoris , en fitta och en ful man , och det var i ett och samma mail .
man behöver inte en doktorsgrad för att se att det lämnar kvar 4 procent för resten av mångfalden .
Japan är världens äldsta land vad gäller snittålder .
det stör mig eftersom jag varit öppen med min homosexualitet ganska länge nu .
och för ett par år sedan bestämde jag mig för att skriva om prokrastinering .
han bestämde att meningen med hans upplevelse var att få känna glädjen i vänskap och sedan lära sig att få vänner .
och jag släpptes .
Hurra ! ni är grymma !
jag hade ett konsultjobb tillsammans med en kollega och vi är så olika som två människor kan vara .
och under nästa decennium kommer vi att ha ytterligare en miljard spelare som är extremt bra på vad det nu än är .
det kan bli otroligt farligt när historier skrivs om eller ignoreras , för när vi förnekas vår identitet blir vi osynliga .
deras konkurrenter är lika kvalificerade att göra alla dessa produkter .
Okej då , vad tror vi om det ?
Vattnet blev hela min värld , varje krusning , virvel , näckrosblad och ström ,
tittar du för mycket på X Factor så köper du kanske idén om att alla kan bli vadhelst de än vill bli .
jag vet inte hur Wagner lyckades med det .
det kan du inte förvänta dig &quot; .
en av 20 personer röstade på vår kandidat som borgmästare i London .
Sperma som finns i kroppen i en vecka eller längre börjar utveckla avvikelser som gör att de inte är lika effektiva på att headbanga sig in i ägget .
vi går tredje året på high school nu , och vi är mentorer åt yngre kårmedlemmar , som en enda sammanhållen grupp .
detta är från Seattle .
vi kan lära oss genom att iaktta andra människor och kopiera eller imitera vad de kan göra .
av respekt för de som kom innan en . gå så här , tala så där , på grund av det .
jag har skrivit en hel bok om det . så jag lever för att lyssna .
Mumier är en fantastisk källa till information , men tyvärr är de geografiskt begränsade och begränsade i historisk tid också .
varför inte ha den snabbtänkthet som Ken Jennings har , särskilt om man kan öka den med hjälp av nästa generations Watson @-@ maskin ?
var så goda och delta i en tyst minut med mig .
jag var orolig för dig när du sa att jag aldrig skulle lämna en tändsticksask någonstans i huset för att mössen kunde komma åt dem och starta en eld .
( musik ) med era 2000 @-@ talsöron föredrar ni det sista ackordet , men förr i tiden skulle ni ha varit förbryllade , irriterade , och några av er skulle ha flytt rummet .
men speciellt i USA väljer många unga bort att skaffa barn och det av samma anledning : ekonomisk oro .
jag samlade pengar i Australien och återvände nästa år för att frivilligjobba på barnhemmet i några månader .
och jag tror att det är högst osannolikt att de var långt från amerikanernas minne när de gick för att rösta i november 2008 .
det var en lögn , men det var min verklighet , precis som de bakåtsimmande fiskarna i lilla Dorothys sinne .
men vi envisas med att förväxla objektivitet och subjektivitet som egenskaper hos verkligheten och objektivitet och subjektivitet som egenskaper hos påståenden .
de lärde oss hur man ger mediciner till möss .
först gick det riktigt bra .
Svaret är , givetvis , att om man spenderar 125 miljarder eller 130 miljarder dollar per år i ett land , bjuder man in nästan alla ,
men underliggande makt är inte alls makt .
och oavsett kultur , oavsett utbildning eller annat , verkar de här sju faktorerna vara närvarande när en person är i flow .
jag är fortfarande exalterad över tekniken men jag tror , och jag är här för att lägga fram min teori att vi låter tekniken ta oss i en riktning , som vi egentligen inte vill .
och det är bara fallet lån .
och jag då ?
och den har utvecklats under tiden .
ska vi vara oroliga ?
och på Stanford har man gjort sådan forskning i fem år nu för att dokumentera hur spelande med en idealiserad avatar förändrar hur vi tänker och agerar i verkliga livet , hur det gör oss modigare , ambitiösare och mer målinriktade .
Naturligtvis nyfikenheten , vetenskapsdelen av det . det var allting . det var äventyr , det var nyfikenhet . det var fantasi .
och ja , vi behöver hopp , det är klart vi gör .
är de inte starkare ?
och 100 företag utanför Idealab och försökte att komma fram till något vetenskapligt .
jag överlevde på endast vatten .
vi samlar blod från dem .
de är några av de minsta satelliter som någonsin avfyrats från världens största satellit .
hur förändrar vi transportvägarna - för varor och människor ?
vi har två väldigt tävlingsinriktade , datakunniga företag .
det är en invecklad dans i 28.000 km / h mellan vår kapsel , som är lik en pytteliten bil , och rymdstationen , som är stor som en fotbollsplan .
många av oss går genom livet och försöker göra vårt bästa i allt vi gör oavsett om det gäller arbetet , familjen , skolan eller något annat .
( Applåder ) jag har utlovats förändring sedan jag var barn .
det var mycket svårt , ska du veta , att göra min auktoritet gällande .
om vi stabiliserar sömnen hos de individer som ligger i riskzonen så kan vi helt säkert göra dem friskare men också lindra vissa av de förskräckliga symptomen hos mentala sjukdomar .
för ur den urbana förstörelsen i Port @-@ au @-@ Prince kom en storm av SMS , människors rop på hjälp , bönfallandes för vårt stöd , delandes information , erbjudandes hjälp , letandes efter deras nära och kära .
var jag än kom , kände det som att min fantasi , var den enda resväska jag kunde ta med mig .
deras biblar har en liten inskription , det står &quot; USA:s armé &quot; på dem .
och jag antar att du injicerar det kanske i ett strutsägg , eller något sådant . och sedan väntar du och , hör och häpna , ut poppar en liten dinosaurieunge .
Gatorna översvämmades men folk ville inte missa chansen att delta vid en sådan nationaldag .
( Skratt ) varför framhärdar vi med att göra samma sak om igen och ändå förvänta oss olika resultat ?
Briljant !
när uppgifterna kom tillbaka räknade jag ut betyg .
när detta gjordes - jag ber om ursäkt - jag kommer använda en förlegad jämförelse mellan uppslagsverk och Wikipedia , men jag gör det för att peka på att när vi gjorde denna inventering , var vi tvungna att titta på massiva mängder information .
och i allra första början är inte alls så många berörda. och då får den klassiska sigmodala , eller S @-@ formade , kurvan .
så det är detta som används .
så att fly från det verkliga samtalet kan ha betydelse eftersom det äventyrar vår förmåga till reflektion .
en tredjedel av alla frukter som vi äter är ett resultat av att insekter tar hand om växternas reproduktion .
de kommer behövas för arbete med avancerade skattefrågor och avgörande stämningar .
men det finns en art i Everglades som du , vem du än är , inte kan låta bli att älska , och det är rosenskedstorken .
varje dag bygger alla vi här gudar som har blivit alldeles vildvuxna , och det är dags att vi börjar slå ner dem och glömma deras namn .
Väck dina åhörares nyfikenhet .
under en lång tid har människor sett vetenskap och humaniora som åtskilda .
vilket jag tycker var en intressant idé , teori .
och detta , så klart , är grundvalen i mycket av den österländska filosofin. samt att det inte finns något oberoende själv , skild från andra mänskliga varelser , som inspekterar världen , inspekterar andra människor .
tio år senare , en annan historia : Iranska revolutionen 1979 .
Nuförtiden får ett av 88 barn diagnosen autism , och frågan är varför kurvan ser ut på detta sätt ?
vi gör detta genom att tänka igenom veckan innan vi befinner oss i den .
där , Mina damer och herrar , utvecklas den amerikanska demokratin under Thomas Jeffersons hand .
Okej , så vad är synestesi ?
( Skratt ) desto smalare jag blev , desto längre kunde jag hålla andan .
om civilbefolkningen dödas , om vapnen tar sikte på samhällen kommer det att föda en ond cirkel av krig , konflikt , trauma och radikalisering och den onda cirkeln är mittpunkten av så många säkerhetsutmaningar som vi står inför idag .
( skatt ) så för att ta tag i problemet samlade jag en grupp internationella forskare i Schweiz , Danmark och Storbritannien
idag tycker jag datorer gör motsatsen .
jag skapar bilderna genom att välja bland korten i ett massivt arkiv från satellitföretaget digital Globe .
håll upp den .
jag har identifierat mig på olika sätt - som bisexuell , som lesbisk - men för mig innefattar queer alla lager av den jag är och hur jag har älskat .
vi var ense om att adresser är dåliga .
min etik för att iaktta är formad av 25 års erfarenhet av att rapportera om tillväxtekonomier och internationella relationer .
och när jag säger &quot; väldigt vanligt &quot; kan det fortfarande vara så sällsynt att inte en enda ö av liv någonsin möter en annan , vilket är en sorglig tanke .
så den kvällen , la jag ut det på Facebook och frågade några av dem , och på morgonen hade svaret varit så överväldigande och positivt , att jag visste att jag måste prova .
Syntetisk biologi , till exempel , strävar efter att beskriva biologi som ett designproblem .
vi måste omdefiniera i grunden vilka som är experter .
hon var dotter till människor som faktiskt varit slavar .
det hade pH 11 , och ändå levde kemosyntetiska bakterier i det . i denna extrema miljö .
vi är inte färdiga med videon än .
när du rör din arm så här , skickar hjärnan en signal till dina muskler här .
så tänker jag &quot; nej , nej , jag vill inte ta konstgjorda preparat , jag vill bara se växter och - bara visa mig örter och växter . jag vill se alla naturliga ingridienser &quot; .
vissa är mindre .
men duvan , som uppenbarligen aldrig gick i flygskolan , sprattlar till , flop , flop , och landar på ena änden av min balansstång .
det är under sömnen vi återställs och återuppbygger oss själva , och när ett hotfullt buller som det här håller på , säger din kropp , även om du lyckas somna , så säger din kropp till dig : &quot; något hotar mig . det här är farligt &quot; .
Föremålet som formade detta var troligen mellan 30 och 50 meter tvärsöver , vilket grovt sett är storleken på Mackeyauditoriet här .
vilket betyder att du kan skapa mening och bygga identitet och fortfarande vara fullständigt ursinnig .
ni ? OK . först av allt , vilket år var det ?
200 miljarder baspar i veckan .
Psykoanalytisk psykoterapi fyra @-@ fem dagar i veckan i decennier och fortlöpande , samt utmärkt psykofarmaka .
ett svar min fru kunde ha gett .
rättigheterna vinns inte i rättssalar , utan i människors hjärtan och själar .
det skulle bli ett köpcenter , istället för en grön oas .
vi kallar varje avläsning för en emotionell datapunkt , och de kan aktiveras tillsammans för att visa olika känslor .
men en sak jag är riktigt nervös för är Mina skakande händer .
jag växte upp med en mycket berömd farfar , och vi hade en sorts ritual därhemma .
LED @-@ lampan strömmar nu videon genom att ändra dess ljusstyrka på ett subtilt sätt. ett sätt som inte uppfattas med vanlig syn , eftersom förändringarna sker för snabbt för att märkas .
det här slog mig när jag skulle köpa nya jeans .
i Ryssland anses jag vara en gammal nucka som aldrig kommer att bli gift .
och att man inte kan existera i det här universumet utan massa .
Ritualerna var bekanta .
och jag tror att TV:n är som en Global lägereld .
i kvantvärlden behöver du inte kasta den över muren , du kan kasta den mot muren , och det finns en viss icke @-@ noll sannolikhet att den försvinner på din sida och dyker upp på den andra .
ta , till exempel , ljudet av ett skott .
vi kommer inte att bryta med dig , och det är något jag alltid har velat att du ska veta , att du är älskad .
det har gett oss motivation till att fortsätta att jobba på detta .
så bara en vecka efter Bergenbanan , ringde vi företaget Hurtigruten och började planera för nästa program .
jag är inte en religiös eller särskilt andlig person , men i vildmarken , tror jag att jag upplevt religionens födelseplats .
( Skratt ) inte för att jag är en dålig lärare , utan för att jag har studerat mänskligt avfall och undervisat i hur avfall transporteras genom reningsverk , och hur vi bygger och designar dessa reningsverk för att skydda ytvatten , till exempel floder .
det var en rätt fantastisk upplevelse , men det är fyra år sedan nu .
när du kombinerar vetenskapen bakom att känna igen bedrägeri men konsten att titta , lyssna , befriar du dig dig från att samarbeta i en lögn .
SM : Ah , ett drag av klassisk övervakningsekonomi .
han bodde i ett område med få vägar där det rådde en stor brist på sjukvårdare .
Extas är alltså att man går in i en alternativ verklighet .
vi kyler ner våra system till nära absoluta nollpunkten , vi utför våra experiment i vaakum , vi försöker isolera dem från alla yttre störningar .
men har vi nått vårt mål ?
vi kan surfa på nätet anonymt .
i stället var det min välsignelse och förbannelse att bokstavligen bli människan i tävlingen mellan människa och maskin som alla fortfarande pratar om .
när vi funderar över konsekvenserna av det och vi tror på att utrotning är vanligt och naturligt normalt och uppstår då och då blir det i högsta grad moraliskt rätt att ha en mänsklig mångfald .
så jag ber er att sprida informationen och håll ögonen öppna .
ett ärligt svar för några månader sedan hade varit , &quot; Vi har ingen aning &quot; .
Thailand , 64 procent .
på Comic @-@ Con eller någon annan Con fotar man inte bara folk som går omkring .
men sedan förstod jag , det är det redan .
Lycka till den här veckan .
jag skulle vilja lägga denna typ av fredagskväll @-@ i @-@ baren @-@ diskussion åt sidan och få dig att faktiskt kliva in i labbet .
Fienden har en röst .
gör som jag , är ni snälla .
2004 så producerade de amerikanska drönarna totalt 71 timmar övervakningsvideo för analys .
Studenterna åkte dit i förväg , och de ordnade så att alla skulle beställa Feynman @-@ smörgåsar .
och dagar har blivit till månader , månader till år .
jag fick lämna dem utan ett ordentligt avsked .
&quot; Oh förlåt , jag blev lite sen . hur går det ? &quot;
Äktenskapsmäklaren tänkte igenom allt , sammanförde två personer , och så var det bra med det .
jag säger &quot; Gud , jag önskar verkligen att jag hade kopplat ihop John Locke &apos; s teori om äganderätt med de efterföljande filosoferna &quot;
om vad ?
och du borde ha alla nätverk från alla dessa relationer mellan dessa element av data .
och nu har vi många bakteriestammar i vår frysbox som får koraller att gå genom den där bosättningsprocessen .
vi reste till byn för att mobilisera samhället .
min fru började bötfälla mig på en dollar för varje irrelevant fakta jag förde in i vår konversation .
eleven försökte , lyckades nästan , men fick det inte att bli alldeles korrekt .
och du har inte varit dig själv .
Landskapet har sorgligt nog befolkats med fler fall som mitt , oavsett om någon har gjort ett misstag eller inte , och nu berör det både offentliga personer och privatpersoner .
att bli blind satte dem i fokus .
Ryan Holladay : Blanda utan skarvar .
och det kanske låg lite sanning i det där , för jag trodde att om jag bara började gå så skulle alla andra , ni vet , följa med .
i filmer är det helt annorlunda .
( Skratt ) och sedan odlade vi celler på dem .
du kan alltså ha inte bara &quot; bilceller &quot; , utan &quot; Aston Martinceller &quot;
mitt sätt behöver dem inte .
människorna .
( musik ) God eftermiddag .
men mycket viktigare , fördelningen är mycket bredare .
redan som barn förstod jag vilka förväntningar som fanns på mig .
jag var inte för juridik .
den har allt inbyggt , och den hoppade för att en student tände en bordslampa bredvid den .
de kommer att vara tillgängliga via maskinen .
Datan visade att jakten på lycka kan göra människor olyckliga .
så därför . om du ser här , nu kan jag fortfarande se det .
de jämförde Dreyfus handstil med den på anteckningen och drog slutsatsen att de stämde överens , även om professionella handstilsexperter utanför det militära var mycket mindre övertygade om likheten , men strunt i det .
KKM : jag har tvingats påminna mig om en massa saker , jag också .
vi behöver tusentals åklagare för att se detta och skydda dem .
men om vi kan få den data ut från bakom fördämningen så att mjukvarutvecklare kan hoppa på dem , på det sätt som dessa utvecklare gillar att göra , vem vet vad vi då kommer att få fram .
mitt favoritexemple är en borrmaskin . vilka här äger en borr , en hemmaborrmaskin ?
vi fick veta att han hade en lång bakgrund av våld i hemmet .
Missförstå mig inte , det vore jättehäftigt att hitta utomjordingar .
här fattas just nu beslutet att du förmodligen inte kommer beställa stek till middagen .
det är ett praktexempel på vad som händer när regeringar attackerar deras egna medborgare . DigiNotar är en certifikatutfärdare
Tyvärr är det inte slutet på historien .
( Skratt ) ca : Sa han att du skulle hoppa , eller var det mer som &quot; jag drar nu !
de är faktiskt skadliga .
och du log mot den jävla kameran som de sa till dig att göra eller så kunde du kan säga hejdå till din födelsedagfest . men ändå , jag har en enorm stapel
det finns människor - några har jag redan nämnt - som är fantastiska , som tror på kvinnors rättigheter i Saudiarabien , som försöker och som får ta mycket hat eftersom dom tar ton och gör sig hörda .
men det finns 22 länder där man talar arabiska och de använder modern standardarabiska , som är den arabiska som används i hela regionen i tidningar och i TV och radio , men självklart skiljer det sig åt mellan länderna i vardagsspråket i dialekter , vardagsuttryck , och så vidare .
vi kan kalla honom Miguel . hans namn är faktiskt Miguel .
( jag är hungrig ! )
de får dig att betala mer i källskatt bara för att bättra på deras pengaflöde .
här är ett foto på mig - jag är överlycklig .
icke @-@ statliga organisationer förstår fördelarna med att ha reportar som följer deras arbete vid sidan om .
Trappistmunken Thomas Merton frågade under Apolloperioden , &quot; Vad kan vi vinna på att segla till månen om vi inte förmår korsa avgrunden som skiljer oss från oss själva ? &quot;
vi behöver transformerande förändring .
den klimatrelaterade extrema torkan som började 2006 i Syrien ödelade 60 procent av jordbruken i Syrien , dödade 80 procent av all boskap , och tvingade 1,5 miljoner klimatflyktingar till Syriens städer , där de kolliderade med ytterligare 1,5 miljoner flyktingar från Irakkriget .
för att lyckas behöver vi alla tillsammans hjälpa och påverka våra politiker , eftersom utan långtgående , världsomspännande förändring så kommer det inte att hända något .
Istället säger de . &apos; nej , nej nej !
i Bangladesh finns ett område som heter Matlab .
året efter , 1949 , gjorde vi beslutet permanent i den nya författningen , och det är därför jag kan berätta denna historia nästan 70 år senare .
( Skratt ) just nu har vi väldigt lovande pilotdata .
vi använder förstås elektricitet . men vi har en lösning åt er - Vi använder oss av en ren energikälla .
2000 år senare kan vi förklara vad som händer i hjärnan .
om vi gör så här tillräckligt ofta , och vi gör det med respekt , kommer folk att tänka efter lite mer kring hur de sätter ihop mötesinbjudningar .
jag frågade dem varför .
en gång tvittrade jag , var i Lembourne kan jag köpa en netiflaska ?
det här är EMMA Ott .
och vi kommer bara att bli tio miljarder i världen , om de fattigaste människorna kommer ur fattigdom , att deras barn överlever och att de får tillgång till familjeplanering .
Istället för att arbeta i samklang med min omgivning , motarbetade jag den .
en garderob är bara ett svårt samtal och även om våra ämnen varierar oerhört mycket , så är upplevelsen av att vara i , och komma ut ur garderoben , universell .
det var en plåga .
så tänk om jag istället för att låta folk summera enskilda TEDTalks till sex ord , gav dem 10 TEDTalks på en gång och sade , &quot; Sammanfatta dessa med sex ord åt mig &quot; .
snart , hoppas vi , ska Masa få återförenas med honom i Sverige , tills dess tas hon om hand på ett vackert barnhem i Aten .
det är faktiskt så att antalet människor som är inblandade i att tillverka en bil har ändrats ytterst lite de senaste årtiondena , trots robotar och automation .
Donald gav oss några av dessa läxor .
skulle vi använda vår auktoritet och makt för att försöka kontrollera eleverna för att hindra dem från att gå , eller skulle vi stötta dem då de utövade de principer om social rättvisa som vi undervisat om sedan årskurs 9 ?
och en av dem är att jag klarar mig bra .
men det är en enorm skillnad mellan Afghanistan och Sri Lanka .
Okej , så ni förstår tanken .
kan det stämma ? det gör det . han var 33 , 38 och 63 när de gjordes .
och den här tävlingsretoriken är standard nu .
men man kan bygga ett godtyckligt antal tunnlar , hur många nivåer som helst .
och sedan byggde hon huset .
för jag vet inte om det finns något värre när det gäller den globala folkhälsan än att låta barn på denna planet dö av sjukdomar som kan förebyggas med vaccin , vaccin som kostar en dollar .
så vi vet att de här kråkorna är riktigt smarta , men ju mer jag grävde i det här , ju mer upptäckte jag att de har gjort en till och med ännu viktigare anpassning .
Låt mig gå igenom dessa tre saker .
män drabbas av autism fyra gånger oftare än kvinnor och vi kan verkligen inte förstå vad som orsakar detta .
de tappade lusten långt innan de har kommit hit .
jag minns att Mina sköterskor klagade på att köra genom det .
Spejaren är den som går ut , kartlägger terrängen och identifierar potentiella hinder .
varför designar jag inte något som mäter fuktnivån i såret så det kan hjälpa läkare och patienter att behandla såren bättre ?
även om vi kunde mäta vad varje cell gör i varje givet ögonblick , måste vi fortfarande få ordning på mönstret i den inspelade aktiviteten , och det är så svårt , risken är att vi kommer förstå precis lika lite av dessa mönster som hjärnan som producerar dem .
vi ska göra detta på människor som har kognitiva störningar och vi valde att behandla patienter med Alzheimers som har kognitiva brister och minnesförlust .
de försvinner på grund av att vissa företag inom skogssektorn går in och skövlar allt .
det var det vanligaste svaret som vi fick .
och istället för att använda magneter eller muskler för att få den att röra sig så använder vi raketer .
Leopardsälen har sedan Shackletons tid haft dåligt rykte .
när jag studerade i Italien , insåg jag att jag saknade arabiskan .
och i en bakterie gör CRISPR @-@ systemet det möjligt att plocka ut DNA:t från viruset och integrerat i små bitar in i kromosomen - i bakteriens DNA .
den ena är att de är mycket vanliga .
så två saker i det här slog djup an hos mig .
nummer ett : vi måste börja göra våldsbekämpningen till en självklarhet i Kampen mot fattigdom .
och deras ledare , deras ledare : innan de skickar sina söner och döttrar att kriga i ert land - och ni vet varför - innan de skickar iväg dem går de till en kristen kyrka och ber till sin kristna gud och ber om skydd och vägledning från den guden .
de föddes alla in i den eller så har de aktivt strävat efter att omge sig med rätt folk .
så medlemmar i mitt team reste omedelbart ut och anslöt till Dr. Humarr Kahn och hans team , och vi möjliggjorde för diagnostisering med känsliga molekylära tester för att fånga upp ebola vid gränsen in till Sierra Leone .
att acceptera det faktum att vi är djur får en del potentiellt skrämmande konsekvenser .
om man tar någon som Portia de Rossi , till exempel , så är alla överens om att Portia de Rossi är en mycket vacker kvinna .
Räck upp en hand om du är i 20 @-@ årsåldern .
det var så , kreativiteten måste hitta sitt utlopp på något sätt .
ute i världsrymden har vi nu en människotillverkad sattelit , som uppenbarligen sänder ut någon slags signal . om vi hittar rätt våglängd kan vi nog höra den &quot; .
jag började ta fram en ny typ av fjärrstyrning . med robotars hjälp kunde jag vara på flera ställen samtidigt- -utan att behöva ta mig dit själv .
Notera bokens titel , &quot; Boken som aldrig checkades ut : Titanic &quot; .
( skratt ) jag tänkte &quot; ja , det är fantastiskt , för jag känner mig inte handikappad &quot; .
jag blev tvungen att leva med två helt olika bilder av mig själv som person ; som en skurk hemma i mitt hemland och som en hjältinna i världen utanför .
när Patrick kom ut från fängelset hade han en olidlig resa framför sig .
jag har investerat i Pakistan i över sju år nu , och de av er som också arbetat där kan skriva under på att pakistanier är en otroligt hårt arbetande folk , och det finns ett häftigt avancemang uppåt i deras natur .
i vårt land . för ytterligare bevis kan vi se på fängelsestatistik ; vi kan se på statistiken över polisvåld gentemot svarta ; vi kan se på utbildningsklyftan - så ja , social rättvisa hör hemma i skolan .
30 färdigheter kunde rädda 30 miljoner liv före år 2030 .
Krigets framtid innehåller också en ny typ av krigare , och det håller faktiskt på att omdana upplevelsen av att gå i krig .
vi har än så länge inga genetiskt förändrade människor , men det är inte science fiction längre .
som vanligt talade vi om världsproblemen .
och mitt absoluta favoritord inom denna kategori är &quot; multi @-@ slacking &quot; .
hon har faktiskt en Harvardpsykolog och har behandlats för bland annat affektiv sjukdom
man behöver inte gå till apoteket längre .
om vi nu vill undersöka detta närmare ?
det sista landet - det sista landet i världen som avskaffade slaveri är samma land som jag föddes i , Brasilien .
varför kände jag mig så berättigad att döma henne ?
jag behöver vila den här veckan &quot; , eller &quot; jag behöver crossträna .
Alldeles strax kommer ni höra ett tåg som de inte reagerar på .
det fanns inga incitament för någon att förbättra produkten , eftersom den finansierades av gåvor .
och det är möjligen de största som någonsin hittats .
så när jag tänker vad som är det fundamentala värdet av ett företag som Tesla , skulle jag säga , förhoppningsvis , om den påskyndade processen med ett decennium , möjligen mer än ett decennium skulle det vara en väldigt bra grej .
så vi måste ställas inför denna fråga : hur får vi våra 1900 @-@ talslagar för krig , som är så åldersstigna nu att de har rätt till äldrevård , att hinna ikapp denna teknik från 2000 @-@ talet ?
vi vet till exempel , från forskning , vad som är viktigast för de som är nära döden : komfort ; att känna lättnad , att inte vara en börda för sina kära ; existentiell frid , och en känsla av förundran och andlighet .
se bara på de här vackra , fascinerande varelserna .
ni förstår vikten av det ?
och ni användare ; det gäller oss alla - vi kan kräva teknik som fungerar på det här sättet .
men , jag hoppas att ni håller med mig om att dessa saker som jag precis beskrivit för er , var och en av dem , förtjänar någon form av pris . ( Skratt ) och det är vad de fick , alla fick ett Ig Nobelpris .
Brutus är Venus granne och &quot; ställa till med bråk &quot; är det som hände dagen efter Venus man hade dött , när Brutus bara kom och slängde ut Venus och hennes barn från huset , stal deras mark , och rånade deras marknadsstånd .
mitt dysfunktionella själv kunde faktiskt koppla in till ett annan själv , inte mitt eget . och det kändes så bra .
med åren har verktyg blivit mer och mer specialiserade .
där finns inga stora gravkammare som de flesta kyrkogårdar kräver bara för att formgivningen ska bli lättare för dem .
Jorden kan sedan användas till att skapa nytt liv .
jag vet inte &quot; . ni vet vad det innebär .
dina minnen och associationer och så vidare .
( Skratt ) Arton minuter , uppenbarligen omöjligt .
den till höger är den som får vindruvor .
du verkar tröttna Bob , men håll ut , för här är den verkliga superegenskapen .
och om vi inte lägger tid och uppmärksamhet på det och tillgodogör oss det lärandet och applicerar det på resten av livet , då är det meningslöst .
men de tävlar även efter att de parat sig , med sin sperma .
detta visade sig vara mycket värdefullt 20 år senare då Michael Bloomberg bad mig bli hans stadsbyggnadschef och gav mig ansvaret att omforma hela staden New York .
min &quot; Svart kille &quot; -grej är så bred och så djup att jag i princip kan sortera och lista ut vem den svarta killen är , och han var min svarta kille .
de är som biologiska fönster som lyser och berättar att cellen nyss var aktiv .
allt började i vårt garage .
här är hon , en Hollywoodkunglighet . jag är en tuff unge från Detroit , &#91; Dolly &#93; är en sydstatsunge från en fattig stad i Tennessee , och vi fann att vi var så synkade som kvinnor , och vi måste ha - vi skrattade - vi måste ha lagt till åtminstone ett årtionde på våra liv .
jag kunde rita . jag kunde måla .
och jag tror att när du söker efter ledarskap , måste du se inåt och mobilisera ditt eget samhälle för att skapa förhållanden som öppnar för en ny sorts lösning .
den värms upp under cirka 30 minuter , kyler ned på ungefär en timme .
Dopaminet som strömmar runt när du är positiv , har två funktioner . det gör dig inte bara lyckligare ,
dessa bilder från American Society for Microbiology visar oss processen .
den första är floden av data som skapas av drönare .
som någon som är ganska nära världsrekordet i antal timmar som tillbringats under en magnetkamera kan jag berätta att en förmåga som är väldigt viktig inom MRT @-@ forskning är kontroll över blåsan .
jag deltog i ett seminarium i år med en skådespelande lärare , Judith Weston .
och det andra alternativet som kan bli klart i tid är hushålls @-@ solel kompletterat med naturgas , vilket vi kan använda i dag , kontra batterierna som fortfarande är under utveckling .
&quot; har du nånsin träffat nån som vaknat på morgonen - ( Skratt ) och blivit svart ? &quot;
Tanken var -- med samma utgångpunkt , ett splittrat land -- att samla tecknare från alla läger och låta dem skapa något tillsammans .
så det är bra , men naturligtvis skulle vi ännu hellre hitta ett sätt att påverka funktionen i hjärnregionen , och se om vi kan ändra på människors moraliska omdömen .
detta var bakslaget i Kenya och Ghana gick förbi , men sedan dalar Kenya och Ghana tillsammans . fortfarande stillestånd i Kongo .
det finns fler : habitatförlust är en av sakerna jag ofta bryter ihop inför mitt i natten .
för mig är de pillren analogin till bilstolarna .
hon säger att det inte finns något mer sinnligt än en het dusch , att varje vattendroppe är en välsignelse för sinnena .
