Om du ansöker om pension från utlandet, får du råd vid Pensionsskyddscentralen.
Kontaktuppgifter till skattebyråns andra serviceställen och telefonrådgivning hittar du på Skatteförvaltningens (verohallinto) webbplats.
Om du vill ha ett arbetsintyg ska du be om det.
Om föräldrarna har ett kombinerat efternamn, blir detta även barnets efternamn.
Skaffa det europeiska sjukvårdskortet i ditt hemland innan du kommer till Finland.
Mer information och råd får du från föreningen Kaapatut Lapset ry.
Att fråga om tillstånd hos hyresvärden om du vill göra ändringar i bostaden, till exempel måla en vägg.
Du får också råd om utarbetandet av en affärsverksamhetsplan och stöd för ditt beslut att starta ett företag.
Om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när hälsostationen öppnar.
Till exempel Sato, Vvo och Avara äger hyresbostäder i Helsingfors.
Oftast betalar hyresvärden förmedlingsarvodet.
Eleverna antas till gymnasiet utifrån vitsorden på avgångsbetyget från grundskolan.
Tolkningfinska
Du kan ansöka till en tionde klass när du har fått ditt avgångsbetyg från grundskolan.
Du kan även registrera bilen på Internet.
Tyvärr kan vi inte svara på respons som är skriven på andra språk.
Företagande kräver yrkeskunnighet och utbildning. Det är viktigt att du är väl insatt i din bransch och lagarna som gäller företagande.
Du kan även besöka mottagningen vid Kliniken för mental- och missbruksvård på servicetorget i Iso Omena utan tidsbokning måndag till fredag kl. 8.30–10.30 och dessutom måndag till torsdag kl. 13–14.30.
Syftet med den partiella sjukdagpenningen är att du kan fortsätta att arbeta eller att återgå till arbetet trots att du har blivit sjuk.
Barnvaktshjälpfinska _ engelska
Du måste beställa tid vid rådgivningarna.
Seure (Seure) är ett bemanningsbolag som erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Hälsotjänster i Vanda
Om du bor i södra, mellersta eller västra Helsingfors finns hälsocentralsjouren vid Haartmanska sjukhuset.
Ta reda på begränsningarna innan du för in läkemedel i Finland.
Unga i åldern 13–23 med missbruksproblem kan få hjälp vid ungdomsstationen.
personnummer
Kommuninvånarna kan delta i och påverka stadens ärenden vid kommunalvalet som hålls vart fjärde år.
Banken behöver följande uppgifter från dig:
om du ska bo stadigvarande i Finland eller vistas här tillfälligt
Definition av en familj
Giftinformationscentralens telefontjänst är öppen 24 timmar om dygnet.
Med bioavfall avses bl.a.:
Barn vid skilsmässa
Skilsmässa
Den initiala självrisken gäller inte mediciner för personer under 18 år.
krigserfarenheter.
Många organisationer och församlingar bedriver också ungdomsarbete.
Företagsverksamheten startas först när stödet har beviljats.
I Vanda ordnas även många rekryteringsevenemang där arbetsgivarna söker arbetstagare.
Tidsbokningen kan du ringa:
Anmälan utan nätbankskoderfinska _ svenska
Lapplands universitetfinska _ engelska
Gymnasiestudierna siktar till studentexamen (ylioppilastutkinto).
Varken staden eller andra hyresvärdar har skyldighet att erbjuda dig bostad.
Vid hälsostationernas preventivrådgivning (ehkäisyneuvola) får du hjälp med graviditetsprevention och familjeplanering.
Din chef berättar för dig om du behöver ett läkarintyg om sjukdomen direkt eller först från och med den fjärde sjukledighetsdagen.
Våld Problem i äktenskap eller parförhållande
Flerspråkiga biblioteketfinska _ svenska _ engelska
bilda ett kombinerat efternamn av era efternamn.
du är medborgare i ett EU-land, EES-land eller Schweiz och du har
Du kan få kostnadsfri hjälp vid Kyrkans familjerådgivningscentral även på engelska och svenska, även om du inte är medlem i kyrkan.
Teatrar i Esbofinska _ svenska _ engelska
På utbildningsstyrelsens (opetushallitus) webbplats finns en sökmotor med vilken du kan se var och när du kan avlägga examen.
Även minderåriga barn kan boka tid hos läkaren och få ett recept för preventivmedel.
Spara lönekvittona.
Mer information om sport som hobby hittar du på InfoFinlands sida Motion.
linkkiMarthaförbundet:
Tandvårdens tidsbeställning och värkjouren nås vardagar kl. 8–15 på tfn 016 322 2562 eller 016 356 1750. Kvällstid och på veckoslut kan du ta kontakt med läkarmottagningen om du är i brådskande behov av vård.
Vid Grankulla konstskola kan barn och unga studera bildkonst och vid Grankulla musikinstitut kan barn och vuxna studera musik.
Min arbetsgivare hotar mig dessutom med våld.
Äldre människors hälsa, Äldre människor
I Finland anlitar många företag revisionsbyråer.
Partiell förtida ålderspension
Mer information om ledigheterna får du på InfoFinlands sida Familjeledighet.
som en kyrklig vigsel.
Erkännande av examen är avgiftsbelagt.
Processen är mycket snabb och smidig.
Om du bor i höghus eller radhus ska du alltid också komma ihåg att meddela husets disponent (isännöitsijä) att du flyttar.
En demonstration ska anmälas till polisen på förhand.
linkkiFörbundet Utvecklingsstörning:
Fundera noga hur företaget drivs och var och hurdana lokaler företaget har.
Seniorrådgivningenfinska _ svenska
Flyktingstatus får de som beviljas asyl eller som tas till Finland i flyktingkvoten.
Kommunerna
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbete med ett annat uppehållstillstånd
bor permanent i Finland
du är arbetslös eller kommer att bli arbetslös
Tolken ska vara vuxen, egna minderåriga barn kan alltså inte användas som tolk.
Könssjukdomar behandlas i huvudstadsregionen på polikliniken för könssjukdomar i Helsingfors.
Karleby evangelisk-lutherska församlingar erbjuder även hobbyverksamhet för barn och unga, såsom lekparksträffar, klubbar, musikverksamhet och läger.
Avgiftens storlek beror på hur många böcker som är försenade och hur många dagar de är försenade.
Också företagaren har rätt till utkomstskydd för arbetslösa.
Därefter placeras invandrareleverna i en finskspråkig klass i sin närskola.
Du kan också bo hemma och gå på rehabilitering därifrån.
Kandidaten ska vara en person
Om du behöver information om hälsotjänsterna, kan du ringa hälsorådgivningen: (09) 310 100 23.
Vistelsetiden på tre månader räknas alltid från det att du varit utanför Finlands gränser.
Möjligheter att studera det finska eller svenska språket
Arbetarskyddsmyndigheten kan förplikta arbetsgivaren att rätta till brister i arbetssäkerheten som förekommer på arbetsplatsen
Lägg till kontaktuppgifterna till dem.
Förskoleundervisning
Kontakta magistraten på din hemort om meddelandet om rösträtt inte skickas hem till dig.
Observera att listan inte nödvändigtvis innehåller allt som måste göras när du flyttar till Finland.
Fpa:s stöd för boendet är följande:
Som fristående examen (näyttötutkinto) (vuxenstuderande)
Arealen är cirka 240 km2, varav cirka 2 km2 består av vatten.
Gymnasieskolorfinska
Kommunerna tillhandahåller många tjänster för sina invånare.
Enligt lag får man inte beställa läkemedel per post från länder utanför EES-området.
Vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn.
Du får hjälp med jobbsökningen på arbets- och näringsbyrån (Työ- ja elinkeinotoimisto), d.v.s. TE-byrån.
Delta och påverkafinska _ svenska _ engelska
Föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk.
Om du själv bokar tolken och betalar kostnaderna kan du anlita en tolk när som helst.
Skriv ut blanketten på Migrationsverkets webbplats och fyll i den färdigt.
dina rättigheter och skyldigheter
Vem som helst kan ansöka om ett bostadslån hos banken.
Ekonomi- och skuldrådgivningfinska.
I InfoFinland under rubriken Officiellt intyg över språkkunskaper får du information om hur du kan jämföra kursernas nivåer med nivån på den allmänna språkexamen (yleinen kielitutkinto).
Examen vid sidan av arbetet med läroavtal
Verksamhetsställen för handikappservicefinska
Du behöver ändå inte borgensmän för ditt lån om du har sparat ihop en del av bostadens pris på förhand, eller om du har annan egendom som duger som säkerhet för lånet.
Läs mer: När du väntar barn.
Klamydia och gonorré behandlas med antibiotika.
Om du inte är kund hos en mottagningscentral kan du ansöka om stöd hos Migrationsverket.
I de lägre årskurserna har man cirka 20 undervisningstimmar i veckan och antalet ökar i de högre årskurserna.
Dessutom har vissa läroanstalter egna studenthem.
Medborgarinstitut
Information för utländska studerandeengelska
legitimation (till exempel pass)
Öppen ansökan
Hälsovårdscentralen
Du får mer information om rätten till hemkommun på InfoFinlands sida Hemkommun i Finland.
Medier
barn och föräldrar
Teater
ortodoxa kyrkan (ortodoksinen kirkko) eller
Därför skulle det vara bra att barnen hade möjlighet att röra på sig tillräckligt också utanför daghemmet eller skoltiden.
Lagar och avtal i arbetslivet
En utredning om dina språkkunskaper
linkkiJämställdhetsombudsman:
På hälsostationen behandlas de vanligaste psykiska problemen.
KOSEK (Karlebynejdens Utveckling Ab) erbjuder tjänster som nyttar företaget under hela dess livscykel, från och med att starta företagsverksamhet.
I Vanda finns också många andra hyresvärdar, varav de största är VVO, Sato och Avara.
Man kan inte heller föreslå en annan person, till exempel en släkting eller vän, som kvotflykting.
Samtal till huvudhälsostationen styrs till ett och samma telefonnummer, (06) 8287 310.
Adress: Steniusvägen 20, 00320 Helsingfors
de som bor i kollektiv.
Transsexuella personer, transvestiter, intersexuella personer och andra människor med mångfacetterad könsidentitet kan få hjälp av jämställdhetsombudsmannen om de upplever diskriminering.
Stadin ammattiopisto är Finlands största yrkesläroanstalt där man kan utbilda sig inom många olika branscher.
Flyttjänsterfinska _ engelska _ ryska
Hälsostationerna har öppet måndag till fredag kl. 8–16.
Information om anmärkning om betalningsstörningfinska _ svenska _ engelska
Handikappservice och stödåtgärderfinska _ svenska _ engelska
Huruvida du omfattas du av den sociala tryggheten och kan få bidrag påverkas också av om du flyttar till Finland till exempel som
Guiden Välkommen till Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
Om du orsakar skador i bostaden måste du ersätta dem.
Läs mer på InfoFinlands sida Yrkesutbildning.
På stadens webbplats finns information om stadsfullmäktige och dess beslut.
Vård av barn i hemmetfinska _ svenska _ engelska
Information om konsumenträttigheterfinska
yrkesvägledning
Om du söker arbete, bör du anmäla dig till TE-byrån.
Du får närmare uppgifter vid social- och närarbetets verksamhetsställe i ditt bostadsområde (sosiaali- ja lähityön toimipiste).
Appar
Grundskolans övriga stödåtgärder omfattar den övriga stödundervisningen i grundskolan, specialundervisning, individuella studieplaner, flexibel bedömning,
Var kan jag få hjälp?
Information om riksdagenfinska _ svenska _ engelska
Om du är under 16 år och behöver preventivmedel, ta kontakt med hälsovårdaren vid din läroinrättning.
Du får personbeteckningen, när du registrerar dig som invånare hos magistraten.
Diskrimineringsombudsmannens kundtjänstfinska _ svenska _ engelska
Om du har ett tillfälligt uppehållstillstånd (B-tillstånd) som är i kraft kan du få en hemkommun om du kan påvisa att det är din avsikt att bo stadigvarande i Finland.
I lågstadiets högre klasser och på högstadiet får de även välja tillvalsämnen.
Inrikesministeriet beslutar från vilka länder kvotflyktingarna tas.
Om samborna har gemensamma minderåriga barn ska de tillsammans besluta om barnens situation på samma sätt som vid skilsmässa.
Många saker i det finländska samhället förändrades.
Om du inte är säker på huruvida banken ger dig ett lån lönar det sig att gå till banken och förhandla om lånet i god tid innan du köper bostaden.
Du ansöker om visum med en visumansökningsblankett.
I samma lokal finns kundtjänsten Osviitta, där du kan köpa resekort till lokaltrafiken.
I vissa gymnasier ges även mycket undervisning i konstämnen.
Från länder utanför EES-området får du ta med dig till Finland den mängd läkemedel för eget bruk som motsvarar högst tre månaders förbrukning.
Navigatorns Startpunkter erbjuder handledning och rådgivning utan tidsbokning till unga under 30 år.
Webbplatsen asuminen.fifinska _ svenska _ engelska
Studentbostäder hyrs ut av studentbostadsstiftelser, universitetens studentkårer, nationer och vissa andra stiftelser.
Du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv.
Klockan 8.00 betyder prick klockan 8.00, inte klockan 8.10.
Vem kan rösta?
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Enligt Finlands lag är män och kvinnor jämställda.
Du kan göra en anmälan om medborgarskap på internet.
Norrskenfinska _ engelska
Vid skilsmässa kommer man överens om hos vilken förälder barnet har sin officiella adress.
Undervisning i det egna modersmålet för invandrare
Skatteförvaltningen gör en del avdrag automatiskt, men vissa avdrag måste du själv ansöka om.
Om du har det europeiska sjukvårdskortet (European Health Insurance Card, EHIC), behöver du ingen separat försäkring.
Sök till högre yrkeshögskolestudier i den gemensamma ansökan.
Allmänt om fackförbund
Du kan få rehabilitering om ditt handikapp orsakar stora svårigheter att klara av vardagen i hemmet, skolan eller arbetet.
En annan anhörig kan få uppehållstillstånd också om han eller hon levt tillsammans som en familjemedlem till den anhöriga som är bosatt i Finland, innan denna person kom till Finland.
Utbildning för invandrarefinska
Lapplands arbets- och näringsbyrå
Vatten
Till slut anslöts hela Finland år 1809 till Ryssland, efter att Ryssland besegrat Sverige i krig.
Mer information om reglerna i Finland ges av Livsmedelsverket (Ruokavirasto).
Läs mer: Brott.
Läs mer om att grunda ett företag på InfoFinlands sida Att grunda ett företag.
Utbetalningen av semesterpenning baserar sig på kollektivavtalet.
du startar företagsverksamheten först när stödet har beviljats.
För ett bostadslån behövs det vanligen en säkerhet (vakuus).
68300 Kelviå
Ofta kan du utbilda dig på arbetstid och arbetsgivaren kan betala för utbildningen.
vård för att förbättra arbets- och funktionsförmågan
Du kan också göra ditt slutarbete i något företag eller göra en arbetspraktik.
Hjälptelefon: 020 316 116
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
När du ansöker om det första uppehållstillståndet i Finland kan du även be om registrering i det finska befolkningsdatasystemet.
Synskadade
Läs mer på InfoFinlands sida Finska och svenska språket.
Skatteprocenträknarefinska _ svenska _ engelska
Tidpunkten varierar men oftast firas påsk i mars eller april.
Morsdag
Via Wilma kan du ha kontakt med barnets lärare och få information om barnets lärande, prov och frånvaron samt händelser i skolan och om skollov.
Sök en bostad i god tid innan du flyttar till Finland
Arbetsgivaren kan även betala handläggningsavgiften för arbetstagaren.
Barnet får automatiskt finskt medborgarskap vid födseln i följande fall:
I detta fall ska du ansöka om en finsk personbeteckning och meddela din adress till magistraten (maistraatti).
Mer information om personbeteckningen hittar du på InfoFinlands sida Registrering som invånare.
Aktiebolaget är den vanligaste företagsformen i Finland.
Bröstcancerundersökningen görs för kvinnor i åldern 50–69 år ungefär vartannat år och undersökningen för livmoderhalscancer för kvinnor i åldern 30–60 år med fem års mellanrum.
Kontrollera vilket alternativ som är förmånligast för dig.
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I detta fall måste du göra en underrättelse om rörlighet till Migrationsverket.
Bland annat hos bostadsförmedlingen, på internet och i lokala tidningar finns annonser om bostäder som är till salu.
Utländska medborgare
Finlands kulturhistoria kan du bekanta dig med bland annat i Finlands nationalmuseum som ligger i Helsingfors.
Läs mer: Teater och film.
Den kostnadsfria rådgivningen ges på finska och engelska.
Ungdomar kan diskutera frågor kring sexuell hälsa med hälsovårdaren vid sin egen skola.
I Helsingfors finns gott om cykelvägar.
Ubildning vid öppna universitetet i Vandafinska _ svenska _ engelska
På Navigatorn kan någon i personalen hjälpa dig att reda ut saker och ting.
Lägenhetshyrorna är vanligen i genomsnitt 100 euro per dygn.
Därtill utbetalas barnbidrag (lapsilisä) till barnets vårdnadshavare fram till dess att barnet fyller 17 år.
Du hittar anvisningar och mer information om ansökan om uppehållstillstånd för uppstartsföretagare på Migrationsverkets och Business Finlands webbplatser.
Asylsamtalet (turvapaikkapuhuttelu) är den viktigaste händelsen under behandlingen av din ansökan.
Till exempel befinner sig en studerande vars enda orsak till vistelsen i landet är studierna tillfälligt i Finland.
Kommunernas idrottsplatser får användas av alla invånare.
På InfoFinlands sida Var hittar jag jobb? finns information om hur du kan hitta ett jobb i Finland.
Dessutom kan du få stöd, rådgivning och handledning.
Läs mer på InfoFinlands sida Barns och ungas problem.
Karlebynejdens institut, som ägs och drivs av Karleby stad, är ett tvåspråkigt (finska och svenska) medborgarinstitut.
Egenvårdsläkemedel (itsehoitolääke) kan köpas utan läkarrecept.
Mer information om makarnas egendom hittar du på InfoFinlands sida Äkta makars rättigheter och skyldigheter.
Rådgivning för och integration av invandrare
Läs mer på InfoFinlands sida Barn vid skilsmässa.
Arbetsgivaren utser för varje arbetsplats en arbetarskyddschef, som bistår arbetsgivaren i samarbetet med anställda och arbetarskyddsmyndigheter.
Om du har anställning i Finland, är det skäl för dig att ansluta dig till en finländsk arbetslöshetskassa.
Om du är studerande kan du söka hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS.
Bibliotekstjänsterfinska _ svenska _ engelska
Läs mer: Yrkeshögskolor, Universitet.
nivåerna B1 och B2: en självständig språkanvändares språkkunskaper (itsenäisen kielenkäyttäjän kielitaito)
Du får då avdragen i efterskott som en skatteåterbäring.
Medlemskapet i panelen binder dig inte till någonting.
Målet är att främja hälsan och välbefinnandet för de blivande föräldrarna och hela familjen och att stöda familjen inför deras nya uppgift som föräldrar och i växelverkan.
Video om arbetstagarens rättigheter i Finlandengelska _ kinesiska _ arabiska _ thai _ hindi
Hyresbostad
Avfallsinsamlingsstationerfinska
På InfoFinlands sida Val och röstning i Finland finns information om vem som kan rösta i kommunaval.
På arbetsplatser och i skolor serveras lunch vanligtvis kl. 11–12.
Vem som helst kan behöva hjälp om livssituationen är påfrestande.
De är fel som ingen känner till.
Centraliserad tidsbokning per telefon: (06) 8287 400
Församlingarfinska _ svenska
Uppsägning av hyresavtal
Se till att det finns tillräckligt många brandvarnare i ditt hem.
Det är bra att skaffa sig en Internetuppkoppling så fort som möjligt efter att du har flyttat till Finland.
På denna sida finns information riktad till kvotflyktingar.
I Helsingfors kan du bli kund hos rådgivningen om du har ett FPA-kort.
Detta innebär att de inte har rätt till FPA:s förmåner.
Fråga mer vid din förläggning.
Du kan också avsluta studierna efter lägre högskoleexamen.
finns information om hur du kan hitta ett jobb i Finland.
Evenemang i Grankullafinska _ svenska _ engelska
Om din hemkommun är Vanda kan du använda kommunens offentliga hälsovårdstjänster.
skattekort och skattenummer samt rådgivning om beskattningen
Om du arbetar vid sidan av studierna är din arbetstid begränsad.
Spara intygen från dina tidigare jobb och studier.
Dessa dagar kan du dela upp på högst fyra perioder.
Läraren bedömer elevernas framsteg i skolan.
Allmän språkexamen, ASE, är ett språktest för vuxna.
Barn som har ett annat modersmål än finska eller svenska kan få modersmålsundervisning.
Vanda erbjuder ungdomar under 20 år gratis preventivmedel.
Webbaserat material
Dagvård i Helsingforsfinska _ svenska _ engelska
Lapplands yrkesinstitut
Trafikfinska _ svenska _ engelska
Information om Migrationsverketfinska _ svenska _ engelska
På finska duar man oftast.
Det är viktigt att du beskriver allt som hänt så exakt som möjligt.
Många städer har rådgivningstjänster för invandrare med rådgivare som specialiserat sig på invandringsfrågor.
Om du bor i en hyresbostad ska du komma ihåg att säga upp din gamla bostad i tid.
Rysktalande klienter: 020 634 4901 (mån.–fre. kl. 10–12 och 13–15)
Läs mer: Trafik.
Det är bra om paret besöker mottagningen tillsammans.
minst tre års arbetserfarenhet från en lämplig bransch
Om man vill fortsätta studierna därefter och avlägga högre yrkeshögskoleexamen, måste man först skaffa sig tre år av arbetserfarenhet från samma område som examen.
Jag måste flytta ut på grund av skilsmässa.
Information om gymnasiestudierfinska _ svenska
De viktigaste verksamhetsformerna består av ungdomsgårdarna, stora ungdomsevenemang, utflykter, internationella utbyten för ungdomsgrupper och sommarkollon för barn.
kursanmälanfinska
Områdeskoordinatorn berättar om hur undervisningen ordnas och hjälper dig i frågor som rör barnets skolgång.
Bostadsrättsbostäderfinska _ svenska _ engelska
Finland för att bo hos en familjemedlem ska du ansöka om registrering av uppehållsrätten för EU-medborgare på grund av familjeband i tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Befolkning
Åldringar
På magistraten utreder man om det är möjligt att registrera en hemkommun (kotikunta)för dig.
Du har rätt att använda arbets- och näringsbyråns tjänster om du har fått kontinuerligt uppehållstillstånd (A) eller permanent uppehållstillstånd (P).
Du kan dra av låneräntan i beskattningen.
Om arbetsavtalet är tidsbundet binder det båda parterna en bestämd tid, om man inte har kommit överens om möjligheten till uppsägning.
På webbplatsen för MIELI Psykisk Hälsa Finland rf (MIELI Suomen Mielenterveys ry) hittar du information om
festivalarbete
Barnet kan även delta i småbarnspedagogik tillsammans med föräldern i lekparker.
P-EU-tillståndsansökan kan även avslås på samma grunder som permanent uppehållstillstånd.
Du behöver följande handlingar:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
LaNuti linkkiLaNuti:
Information om boendefinska _ engelska
Då är tolkningen kostnadsfri för dig.
Skilsmässa och vårdnad om barn
Överväger du att avbryta graviditeten?
Du krävs inte på redogörelse över din utkomst.
linkkiCIMO:
Läs mer: Stöd- och serviceboende
Det finns också caféer där kunderna har möjlighet att använda Internet.
Nationalparkerfinska _ svenska _ engelska _ ryska _ kinesiska
sexuell läggning.
I början av CV:t kan du tillfoga en sammanfattning eller profil där du beskriver din bakgrund och din kärnkompetens med några ord.
Finskans grammatikengelska
På den här sidan finns information om tjänsterna i Rovaniemi.
Chatbot-tjänst för utländska företagarefinska _ engelska
Påsk
Bästa stället att fråga om enskilda grenar och var man kan utöva dem är grenförbunden.
Ta med dig identitetsbevis och uppehållstillstånd.
Sporrgränden 2 A, vån. 3 (Håkansböle)
Du kan också vända dig till Huvudstadens Skyddshem (Pääkaupungin Turvakoti).
FPA ordnar rehabiliteringen och ersätter kostnaderna för den.
Privat psykoterapitjänst på Internetfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ norska
En brandvarnare kan rädda ditt liv.
Barn kan också gå i en skola med en speciell inriktning.
Hen ger dig råd och ser till att dina rättigheter förverkligas.
När en person som är fast bosatt i Finland blir arbetslös, har han eller hon rätt att få utkomstskydd för arbetslösa.
Förmånligast övernattar man i delat rum.
Bostäderna är dyrare nära stadens centrum.
Om man bryter mot trafikreglerna kan man få böter.
Finland accepterade resedokumentfinska _ svenska _ engelska
Arbetsgivaren kan ansöka om stöd för arbetstagarnas finskundervisning via arbets- och näringslivstjänsterna.
Skyddshemmet Mona är endast avsett för invandrarkvinnor och deras barn.
De offentliga tjänsterna började utvecklas och på så sätt skapade man den offentliga hälsovården, sociala tryggheten och grundskolan.
För att kunna ansöka om ett nytt uppehållstillstånd för arbetstagare måste du ha ett nytt jobb.
Kindpussar är dock ovanliga.
Dixi, Banvägen 11, 2:a vån.
Du kan prata om dina problem med skolans eller läroanstaltens hälsovårdare eller de vuxna vid ungdomsgården.
Om du vill kan du även be någon annan släkting eller en vän att följa med.
En utvecklingsstörd person som behöver vård kan bo i ett familjehem.
Lapplands yrkesinstitut
tfn (09) 8392 3415
På universitet kan man avlägga lägre högskoleexamen på cirka tre år och därefter högre högskoleexamen på cirka två år.
Helsingfors stad ordnar eftermiddagsverksamhet för barn i årskurs 1 och 2 i skolor och lekparker efter skoldagen.
Tfn 029 55 39391
Myndigheterna överväger beviljandet av uppehållstillstånd alltid fall för fall.
Detta kallas för aktiveringsmodellen för arbetslöshetsförsäkringen (työttömyysturvan aktiivimalli).
Du får stanna i Finland om du beviljas asyl eller uppehållstillstånd på någon annan grund.
Du kan lära dig ett nytt yrke eller en ny examensdel.
Regler
Ansvarig bolagsman i kommanditbolag
Finlands utrikespolitik i samverkan med statsrådet och
Grundläggande information om yrkeshögskolorfinska _ svenska
Du har möjlighet att få en hemkommun i Finland om:
Dessa nivåer delas ytterligare in i undernivåer.
Passfoto (anvisningar för fotot finns på Migrationsverkets webbplats)
På hjälptelefonen får du stöd och vid behov råd om var du kan få hjälp.
Konserterfinska _ svenska _ engelska
Privata mentalvårdstjänster
Läs mer: Högskoleutbildning.
Företagsverksamhet som bisyssla lönar det sig ofta att starta som enskild näringsidkare.
Separat insamlat bioavfall packas i en papperspåse, en påse vikt av en dagstidning eller en plastkasse. Kassen eller påsen får vara högst 30l stor.
Invånarhusen Kivenkolo och Kylämaja är öppna för alla.
För dessa koder gäller dock hårdare krav än för öppning av ett bankkonto.
Du kan även söka fram en privat advokat via Finlands Juristförbunds webbplats.
Om bostaden är större eller dyrare än vad lagen om allmänt bostadsbidrag tillåter växer den andel av boendekostnaderna som du betalar själv.
För att teckna ett abonnemang behöver du ett finländskt identitetsnummer och du måste ha en adress i Finland.
På utbildningsstyrelsens (opetushallitus) webbplats finns en sökmotor för språkexamina.
Öppet varje dag dygnet runt.
Bildkonst
Dessutom krävs att:
Ta i god tid reda på när du kan ansöka om en studieplats.
Övriga länders medborgare måste anmäla sig personligen hos TE-byrån.
Då ordnas fyrverkerier.
Kvinnan har rätt att själv besluta om hon vill göra abort.
Då kan domstolen döma till skilsmässa direkt.
Hur ordnas umgänget?
En besvärsanvisning om hur beslutet får överklagas bifogas alltid beslutet.
Läs mer om sjukförsäkringen i Finland på InfoFinlands sida Den sociala tryggheten i Finland.
Utbudet kompletteras av språk- och metodstudier.
I hälsovården av barn under skolåldern får man hjälp av rådgivningsbyråerna (neuvola).
Diskriminering (syrjintä) är ett brott.
På Finlex webbplats kan du läsa lagen angående vårdnad om barn och umgängesrätt.
Studierna omfattar mycket praktiska övningar.
Privat dagvårdfinska
Telefon: 029 56 49294
Vid vårt vetenskaps- och konstuniversitet fås utbildning och idkas forskning inom pedagogik, turism och affärsverksamhet, juridik, konstindustri och samhällsvetenskaper.
Europass är särskilt nyttigt om du ansöker om ett jobb eller en utbildningsplats i Finland från ett annat EU-land.
När du ansluter dig till ett fackförbund kan du samtidigt ansluta dig till förbundets arbetslöshetskassa.
Det finns inga möjligheter att övernatta på nattcaféet, och det är inte heller drogfritt.
Hälsostationernas adresser:
Du kan använda de offentliga hälsovårdstjänsterna om du har en hemkommun i Finland.
På InfoFinlands sida Att grunda ett företag hittar du information om hur man grundar ett företag i Finland.
För hormonella preventivmedel behöver du ett recept av en läkare.
Familjeledigheter
Hälsostationen på Rinteenkulmafinska
Också sökandens inkomster beaktas, eftersom bostäderna främst är avsedda för personer med låga inkomster.
Utbildning som handleder för yrkesutbildning (VALMA)
Samhället tryggar barnets rättigheter med hjälp av lagar och författningar.
Enligt Finlands lag ska alla människor behandlas likvärdigt oberoende av deras bakgrund och kön.
Det åligger kommunerna att ordna serviceboende och stödboende för personer som behöver det.
Du kan ta direkt kontakt med en arbetsplats som du är intresserad av.
Läs mer:
Ibland är dessa skolor privatskolor.
Finska medborgares rättigheter och skyldigheterfinska _ svenska _ engelska
Din uppehållsrätt kan registreras om du är anställd eller har ett eget företag i Finland.
Det har på grund av förälderns ekonomiska situation fastställts att inget underhållsbidrag betalas.
Avtala om arvodet skriftligen på förhand.
Studentexamen består av prov i olika läroämnen.
Du får alltså både yrkesutbildning och en arbetsplats.
Juristens rådgivning per telefon 020 316 117
Diabetes kan behandlas med insulin och rätt kost.
Att röra sig i naturen
Förete skattekortet till din arbetsgivare.
Mer information hittar du på FPA:s webbplats.
Hyresbostäderfinska _ svenska
hör till en finländsk arbetslöshetskassa
Vid Esbo musikinstitut (Espoon musiikkiopisto) kan barn och vuxna studera musik.
du har tidigare haft en hemkommun i Finland
I staden finns flera busslinjer.
De flesta utrikesflygen avgår från Helsingfors-Vanda flygplats.
Läs mer på InfoFinlands sida Dödsfall.
Kasta inte avfallet ut genom fönstret, i skogen eller på gatan.
Du hittar jobbförmedlingssidor när du skriver "avoimet työpaikat" (lediga jobb) i sökmotorns sökfält.
Migrationsverket skickar dig en kallelse till asylsamtal.
De högsta tjänstemännen i Rovaniemi stad är stadsdirektören och två biträdande stadsdirektörer.
I Finland kan du studera på finska, svenska och ibland på engelska.
Sådana preventivmedel är till exempel p-piller och minipiller.
Förskoleundervisningen är avsedd för sexåringar och den ges vid daghem.
När du har en hemkommun kan du använda kommunens tjänster, såsom till exempel hälsovårdstjänster.
ryska och engelska tfn 050 325 7173
Det allmänna nödnumret är 112.
Om du är sambo med en finsk medborgare som bor i Finland kan du få uppehållstillstånd på grund av familjeband.
Du kan även ta dig till Huvudstadens Skyddshem.
Evenemang och sevärt i Helsingforsfinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Söka bostad
Ainonkatu 1, vån.
Enligt lag får ingen diskrimineras till exempel av följande orsaker:
Att ansöka om skilsmässa
Du får mer information om tolktjänsterna i din kommun på rådgivningsbyrån.
Presidentval
Låt göra en läkarundersökning före utgången av den fjärde graviditetsmånaden.
När Migrationsverket har gett ett positivt beslut på din ansökan om återförening på grund av familjeband och anser att staten kan bekosta resan för dina familjemedlemmar, skickar det sitt beslut till Röda Korset.
Observera att tull- och skattefriheten för flyttsaker inte gäller alkohol eller tobaksprodukter.
Motion
Till reglerade yrken hör både uppdrag inom den offentliga sektorn och yrken för vilka det krävs rätt till yrkesutövning.
Du kan studera finska eller svenska.
Då firas i Finland midsommar, som är midnattssolens och högsommarens fest.
En utredning om ditt uppehälle.
På Omnia ordnas för invandrare utbildning som förbereder dem på yrkesutbildning.
Nylands arbets- och näringsbyrå, Esbo
vistas i landet illegalt
I arbetslivet ska kvinnor och män behandlas lika.
Tfn (09) 839 21074 och (09) 839 32042
Vuxna invandrare som inte har grundskolans avgångsbetyg från sitt eget land kan avlägga grundskolan på vuxengymnasiet.
Det kan variera allt mellan dagliga till veckovisa hembesök.
Nollalinja är en hjälptelefon som du kan ringa om du har blivit utsatt för våld i familjen, sexuellt våld eller hot om våld.
Barnskyddslagen (Lastensuojelulaki) säger att alla barn bosatta i Finland har rätt till omsorg och en trygg uppväxtmiljö.
Rehabiliterande psykoterapifinska _ svenska _ engelska
Företagare som säljer varor och tjänster i Finland är skyldiga att betala mervärdesskatt.
Fångstvägen 3
Bio Rex program finns under länken här intill.
Vid yrkeshögskolorna och universiteten i Esbo och Helsingfors kan du studera inom många områden.
rehabiliteringspsykoterapi
Om du blir arbetslös
Studierna på studielinjerna pågår i 1–2 år.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kontakta ett skyddshem.
Människohandelns offer kan få hjälp.
Om du inte korrigerar skattedeklarationen, förblir det här beskattningsbeslutet i kraft.
Om du inte betalar räkningen senast på förfallodagen eller inte har kommit överens om att förlänga betalningstiden, måste du betala påminnelse- och inkassokostnader samt dröjsmålsränta.
Exporten av tjära, som blev mycket viktig för Karlebys historia, inleddes redan på 1500-talet.
Att köpa sexuella tjänster av ett barn under 18 år är ett brott.
Tidsbeställning
Största delen av läkemedelsbutikerna på internet är dock illegala.
Om du har en funktionsnedsättning, ta då först kontakt med hälsostationen (terveysasema).
Velkalinja är Takuusäätiös kostnadsfria rådgivningstelefon.
67701 Karleby
Meddela numret på ditt bankkonto via Skatteförvaltningens webbtjänst eller på en separat pappersblankett.
Intern kommunikation på arbetsplatsen
Av det ser arbetsgivaren, hur mycket skatt som ska betalas på lönen.
Den är gratis.
Finlands förhistoria –1323
På InfoFinlands sida Våld hittar du information om vad du kan göra om din partner utövar våld eller hotar med våld.
Du måste meddela daghemmet och skolan när barnen slutar där.
Mariegatan 16–20 (l-flygeln, ingång B1)
Hyresvärden har hotat med att vräka mig från hyresbostaden på grund av högljutt liv.
Kvällar och helger
Du kan söka till en yrkesutbildning när du har avlagt lärokursen för den grundläggande utbildningen.
Etableringsanmälan
Läs mer: Hyresbostad.
Om din närstående utgör en fara för sig själv eller för andra och inte går med på att träffa en läkare kan du ringa hälstocentralen eller sjukhuset.
Förlossningfinska _ svenska _ engelska
Polikliniken för könssjukdomarfinska _ svenska _ engelska
Om säljaren av bostaden godtar köpeanbudet görs bostadsköpet upp i köparens bank.
Mer information om möjligheter till musikhobby får du via kommunens kulturkontor.
Den internationella föreningen i Håkansböle (Hakunilan kansainvälinen yhdistys) har en rådgivningspunkt som betjänar invandrare i Håkansböle, Björkby och andra områden i Vanda, som vill ha information om till exempel studier, språkkurser, arbete, hobbyverksamhet, krissituationer eller juridiska frågor.
Du kan inte få flexibel eller partiell vårdpenning om du får föräldradagpenning och/eller hemvårdsstöd och själv tar hand om dina barn.
Folket kom österifrån från nuvarande Rysslands område och söderifrån via Baltikum.
Karleby finska gymnasium erbjuder förberedande undervisning för gymnasiet även för invandrare.
omfattas av den finländska sjukförsäkringen (sairausvakuutus): läs mer på InfoFinlands sida Den sociala tryggheten i Finland
Information om finska romanifinska
På daghemmet är barnen i större gruppen är i gruppfamiljedagvården.
Folk flyttar till Finland
Delägare som innehar en ledande ställning i ett aktiebolag (verkställande direktör eller styrelsemedlem) eller person som innehar en ledande ställning i någon annan sammanslutning
Skrapning görs vanligtvis i narkos och därefter ska du stanna några timmar på sjukhuset.
Måste jag betala?
Du kan även fråga om mer information av daghemsföreståndarna.
Minnesstörningar och demensfinska _ svenska _ engelska
Fråga om råd på företagsrådgivningen
dina inkomster inte är för stora; och
FPA
Den närmaste byrån finns i Esbo.
Man kan ansöka om bodelningsman om samboförhållandet har varat minst fem år och parterna har gemensamma barn.
Gymnasiet är en allmänbildande utbildning som inte ger ett yrke.
Publikationer eller andra arbetsprov
Tfn 09 3104 4556 (mån–fre kl. 9–15)
Familjerådgivningscentralenfinska
På stadens webbplats hittar du också anvisningar om hur du söker hyresbostad.
Finskt medborgarskap till barn med finsk farfinska _ svenska _ engelska
Bostadsrättsbostäderfinska
linkkiMetropolia:
Finnkino är den största biografkedjan i Finland.
När du blir sjuk ska du kontakta hälsostationen i ditt område.
Barnkulturcentralen Musikantitfinska _ engelska _ ryska
En studerande från ett land utanför EU/EES kan ha rätt till vissa av FPA:s förmåner, till exempel de förmåner som ingår i sjukförsäkringen.
Hörselapparatfinska
Läs mer: Hälsovårdstjänster i Finland.
Stöd för familjer
Om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen.
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
De ungas skyddshus
I Finland har vi fyra mycket olika årstider.
FPA:s kostnadsersättningfinska _ svenska _ engelska
Ring journumret 045 639 6274 om du behöver en plats på skyddshemmet.
linkkiMellersta Finlands tolkcentral:
Därefter ger TE-byrån ett utlåtande i ärendet till den instans som betalar förmånen, det vill säga till arbetslöshetskassan eller FPA.
Om du vill ha mera kunskap och färdigheter innan du söker till en yrkesinriktad utbildning, kan du ansöka till VALMA-utbildningen.
Också positiva saker, t.ex. att man får barn, kan ändra livet så mycket att man behöver stöd i den nya situationen.
Du kan få stöd för skolresor (koulumatkatuki) om du bor i Finland och studerar i gymnasiet eller vid en yrkesläroanstalt.
Fråga mer vid den läroanstalt där du vill studera.
Patientombudsmannens tjänster är kostnadsfria.
Om du är kund hos en mottagningscentral kan du ansöka om stöd för frivilligt återvändande vid din egen mottagningscentral.
Under samtalet får den som ringer hjälp med att kartlägga sin situation, råd och vid behov vägledning till något ställe där man kan få hjälp.
Rättighet
Som EU-medborgare behöver du inget arbetstillstånd i Finland.
Nybörjarnivån
Kontorets öppettider
Vad kan jag studera i yrkesinriktad arbetskraftsutbildning?
Privat dagvård och hemvårdsstöd
Observera att handlingarna ska vara på finska, svenska eller engelska.
Läs mer: Handikappade personer.
I Finland kan alla gifta sig som
I nödsituationer ringer du det allmänna nödnumret 112.
Du kan fråga vid närmaste FPA-byrå hur du kan få hjälpmedel.
Böcker och annat material finns på flera olika språk.
Om äktenskapet slutar i skilsmässa delas makarnas sammanlagda egendom jämnt mellan makarna.
Fyll i blanketten i Enter Finland-tjänsten.
Brott kan anmälas per telefon eller fax, på polisens webbplats eller genom personligt besök till polisstationen.
Service för missbrukarefinska _ svenska
Arbetsgivaren ska ge den anställda en skriftlig redogörelse för de centrala villkoren i arbetet vid tillsvidare gällande anställningar samt anställningar som varar över en månad.
Du kan resa till Finland om du har ett giltigt ID-kort eller pass.
hittar du en lista över webbsidor där du kan ansöka om bostad.
Uthyrning i andra hand
Läs mer på InfoFinlands sida Universitet.
registrerat uppehållstillstånd;
Läs mer: Trafik.
Rabatter för pensionärer
praktik projekt
Du ska ha med dig kortet på varje besök till rådgivningen.
Socialhandledare 016-322 3124, 040-729 8766
byta en säkring
Fackförbundets representant på arbetsplatsen
Till en del kurser kan du anmäla dig på Internet.
Du kan lära dig ett nytt yrke eller en ny examensdel.
Om en närstående dör oväntat och du behöver stöd kan du kontakta social- och krisjouren i Esbo, telefon (09) 816 42439.
För att barnet ska kunna få uppehållstillstånd måste hans/hennes uppehälle i Finland vara tryggat, till exempel genom förälderns löneinkomster.
Om du redan har finländsk personbeteckning och ett skattekort, hittar du skattenumret på ditt skattekort.
Tfn (09) 505 6379
Företagshälsovårdens tjänster
Den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader.
tillräckliga kunskaper, färdigheter och resurser för den företagsverksamhet som du planerar
Att färdas på isen
Stöd vid skilsmässafinska
Vård av barnet
Teater och filmer
I det här fallet är tolkningen avgiftsfri. Tolkning ska alltid begäras i förväg.
Likväl utreds alla ansökningar som EU-medborgare skickar in.
Läs mer på InfoFinlands sida Diskriminering och rasism.
Du ska då bifoga till ansökan ett löneintyg för löner som du har fått.
Användningen av dem kan vara begränsad, men oftast är de öppna för alla.
Privata hälsovårdstjänster är dock avsevärt dyrare för kunden än offentliga.
Arbetsförmedlingstjänster
Stödboende för personer med psykisk ohälsa och missbruksproblemfinska
Ansökan till förskoleundervisningfinska _ svenska _ engelska
ränteavdrag på bostadslån
på ett daghem (päiväkoti)
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Till exempel får syskon inte ha samma namn som första namn.
CV:t kan även vara en video, en portfölj eller en webbsida.
Enligt lagen i Finland måste arbetstagarna behandlas väl och de ska betalas lön.
Fundera på hur ditt kunnande motsvarar arbetsgivarens önskemål och krav.
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Underhållsbidrag för barn
Bostadssituationen varierar mycket mellan olika orter.
Öppningsoperationen gör förlossningen och undersökningarna under graviditeten lättare.
Du kan läsa mer om registreringen av modern på InfoFinlands sida Registrering som invånare.
Tolktjänster
En meritförteckning, eller ett CV, är en kortfattad och tydlig sammanfattning av ditt kunnande, din arbetserfarenhet och din utbildning.
Vaccinationer är en central del av förebyggandet av smittsamma sjukdomar hos barn. Barnrådgivningen ger barnet de vanliga vaccinationerna.
Sökandens livssituation och behov av understöd är ofta mycket olika.
Du får mer information om tolktjänsterna i din kommun på rådgivningen.
Gör en skriftlig anmälan till din arbetsgivare senast två månader innan du blir moderskapsledig.
Sexuellt våld
Invånarna i Esbo kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
äkta par och registrerade par sambor
Du får arbetslöshetsförmån under utbildningstiden.
linkkiEuropaskolan i Helsingfors:
Giltigt ID-kort eller pass
Läs mer på InfoFinlands sida Uppehållstillstånd för make eller maka.
Rasism (rasismi) innebär att man betraktar någon människogrupp eller en person som hör till gruppen som sämre än andra till exempel på grund av etniskt ursprung, hudfärg, nationalitet, kultur, modersmål eller religion.
Barnen äter tre måltider under dagen: frukost, lunch och mellanmål.
Om barnet inte är tryggt i sitt hem eller om situationen med barnet är mycket svårt, kan det fattas ett beslut om vård utom hemmet eller omhändertagande.
Om du inte har en hemkommun i Finland ska du be FPA utreda din rätt till den offentliga hälso- och sjukvården.
Yrkesubildning
Enkäterna är oftast på engelska, ibland även på andra språk.
Esbo huvudpolisstation
Mer information finns på Karleby kyrkliga samfällighets webbplats.
Arbetsgivaren kan t.ex. betala avgifter för en kurs i finska för din räkning.
Vård av barn Invånarparker och klubbar
Det är bra att inleda medicineringen så tidigt som möjligt.
Läroanstalten meddelar dig att du har antagits för studier med ett brev.
Hörselförbundet och Finlands Dövas Förbund är organisationer som arbetar för att förbättra hörselskadade personers ställning i samhället.
Du får studera i Finland högst 360 dagar när du gör en underrättelse om rörlighet.
Du kan också söka bostad via föreningen Suomen Opiskelija-asunto (Suomen Opiskelija-asunto) (SOA).
Följ väderleksrapporterna och använd alltid en flytväst i rätt storlek.
Du behöver intyget om du ansöker om moderskapsledighet av din arbetsgivare.
Användaren kan förhindra användningen av cookies i sina webbläsarinställningar.
När du har sökt asyl har du rätt att vistas i Finland medan din ansökan behandlas.
Föräldern kan då ha antingen ensam eller gemensam vårdnad om barnet.
Om dina inkomster blir mindre eller större under året, ska du beställa ett nytt skattekort.
Kontrollera regelbundet att brandvarnaren fungerar.
Om du flyttar utomlands för över ett år, betraktas flyttningen som permanent flyttning.
Eldstadsvägen 7 B, vån.
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
Ansökan ska göras innan du har vistats utomlands över två år.
bedömningen av hur bra du kan klara av studierna.
Så här ansöker du om Schengenvisum
Det kallas för lättföretagande.
Möblerade hyresbostäder och lägenhetshotell
yrkesutbildning
via tjänsten Mina e-tjänster eller per telefon.
Arbets- och näringsbyrån anvisar invandrare till kurser i finska språket som ingår i integrationsprocessen.
Socialtjänsterfinska _ svenska _ engelska
Detta innebär att du håller en paus i lyftandet av pensionen.
Mer information om familjeåterförening finns på InfoFinlands sida Till familjemedlem i Finland.
I den inledande kartläggningen får du information om utbildning i finska eller svenska, arbetssökning, utbildning och tjänster i Vanda.
linkkiFöreningen för mental hälsa i Finland:
Ungefär fem procent av finländarna har svenska som modersmål.
Läs mer om finska medborgarnas rättigheter och skyldigheter på InfoFinlands sida Finskt medborgarskap.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Vandainfon finns i Dickursby, Korso och Myrbacka.
Anmälningstiden är i början av året, vanligen i januari.
Grundläggande utbildning
ABC för restaurangbranschen:
I Finland tillhandahåller kommunerna kommunal småbarnspedagogik bland annat i daghem.
När du söker sjukdagpenning ska du bifoga till ansökan:
Hemvårdsstödet består av en vårdpenning och ett vårdtillägg som är beroende av familjens inkomster samt ett eventuellt kommuntillägg.
Människorna samlas på picknick.
Fastställande av faderskap (Isyyden tunnustaminen)
linkkiInstitutet för hälsa och välfärd:
Du kan inte identifiera dig med ett körkort.
Också universitetet flyttades år 1828 från Åbo till Helsingfors.
Kurser – Lista kurserna i finska och andra kurser som du avlagt under en egen rubrik.
I Helsingfors finns det också privata skolor med undervisning på t.ex. engelska, tyska, franska eller ryska.
Från EES-länderna får du ta med dig den mängd läkemedel för eget bruk som motsvarar ett års förbrukning.
Även andra anhöriga till en person som har ett uppehållstillstånd på grund av internationellt skydd kan beviljas uppehållstillstånd.
Förtroendemannen väljs av de anställda.
en hyresbostad
Samtal på finska
Pensionsbeloppet beror på hur länge personen har bott eller arbetat i Finland.
Dit kallas brottsoffret, den brottsmisstänkta och vittnen.
Vissa preparat kan tas inom 120 timmar efter samlaget.
Du kan beviljas asyl i Finland om myndigheterna anser att du blir förföljd i ditt hemland på grund av
utan tvingande skäl göra upp öppen eld på annans mark
Ansökan till vissa universitetsstudier sker genom en separat ansökan.
Dessutom krävs det att du har haft din hemkommun i Finland i minst två år i rad.
Ingen får dömas till döden eller torteras.
En invandrarförening kan hjälpa dig att bevara och utveckla din kultur.
Familjerådgivningfinska _ svenska
Polska
Rättigheter
Umgängesrätten kan till exempel innebära att barnet bor hos den ena föräldern och träffar den andra föräldern vartannat veckoslut och dessutom vissa tider under loven.
Olika konstarter är musik, bildkonst, dans, teater, cirkuskonst, ordkonst, handarbete och arkitektur.
Om du har betalat för mycket i skatt, får du skatteåterbäring (veronpalautus).
Innan du skriver din jobbansökan, läs jobbannonsen noga och fundera på vilka färdigheter och vilket kunnande arbetsgivaren är ute efter.
Den har öppet dygnet runt.
Barn under 15 år behöver ett läkarrecept.
Bybibliotek linkkiBybiblioteken:
Kränkande eller osakligt innehåll
Med hjälp av gränssnittet kan du visa InfoFinlands innehåll på andra webbplatser eller skapa olika applikationer.
Traumatiska upplevelser
Information om tjänsterna finns på sidan Som invandrare i Vanda.
Fredrikinkatu 48
Helsingfors enhet
Hedersrelaterat våld kan vara till exempel
En del områden är väldigt populära. I sådana områden hyrs bostäderna ut mycket snabbt.
Tjänsterna vid A-kliniken i den egna kommunen är kostnadsfria för klienter som bor stadigvarande i Finland.
Regionala ungdomstjänsterfinska
I Helsingfors finns många privata läkarstationer som även tar hand om barn.
du ber en släktning eller vän gå i borgen för ditt lån.
Läs mer om vem som omfattas av den finländska sjukförsäkringen på InfoFinlands sida Den sociala tryggheten i Finland.
Malms sjukhus
Lapplands yrkeshögskolafinska _ engelska
Äldre människors hälsa.
Yrkeshögskolan kan ordna avgiftsfri utbildning för invandrare med målet att ge den studerande tillräckliga språkkunskaper och andra färdigheter som behövs för att studera vid yrkeshögskolan.
På InfoFinlands sida I Finland utan uppehållstillstånd finns det mer information för papperslösa.
Du kan få stöd om du på grund av ditt handikapp eller din sjukdom behöver kontinuerligt hjälp.
Tjänster för handikappadefinska
Privata hyresbostäder
Om du misstänker att ett barn har förgiftats kan du fråga råd vid Giftinformationscentralen (Myrkytystietokeskus).
Företagarens skyldigheter
För akutpreventivmedel behövs vanligen inget recept.
Problem i skolan eller med studierna
På gymnasiet behövs goda språkkunskaper.
Broschyren Att söka pension från utlandetfinska _ svenska _ engelska _ ryska _ estniska
pedagogiska områden
År 1946 inkorporerades nya områden till Helsingfors och staden yta mångfaldigades nästan åtta gånger.
Om du insjuknar plötsligt eller om du råkar ut för en olycka, får du akut sjukvård även om din hemkommun inte är Vanda.
Stämpeln ska begäras vid utrikesministeriet i det ifrågavarande landet och dessutom vid Finlands beskickning i landet.
Du kan ringa brottsofferjouren om du eller en närstående har blivit utsatt för ett brott eller om du har bevittnat ett brott.
Telefonrådgivning: (09) 816 45285
arbetsgivarens och arbetstagarens hemort eller driftställe
Karleby handelsflotta var under perioder Finlands största.
Ekonomi- och skuldrådgivning ordnas av kommuner.
Ett försäkringsintyg eller en kopia av det europeiska sjukvårdskortet
MoniNet är ett mångkulturellt center i Rovaniemi, Lappland.
Rådgivningsbyrån för familjeplanering ger stöd i frågor om familjeplanering och graviditetsprevention.
Stöd till företagare
Du får information om hur du köper läkemedel på InfoFinlands sida Läkemedel.
Arbetsgivaren måste följa kollektivavtalet.
Information om hälsorådgivningfinska _ svenska _ engelska
Rådgivningen betjänar telefonledes på numret 045-237 7104 (måndagar kl. 14–16).
Naturens husfinska _ svenska _ engelska
linkkiVanda stad:
På samma adress ser du också hur behandlingen av din ansökan framskrider.
Om du till exempel orsakar en vattenskada måste du själv betala hela renoveringskostnaden.
I studiemiljön finns sju avsnitt som handlar om invandrarens liv i Finland.
Vilka reklammedel ska du använda för att främja försäljningen?
Rehabiliteringsstöd är invaliditetspension på viss tid.
Läs mer: Fortsatt uppehållstillstånd.
I Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig.
Erkännande (BY) – Du måste nämna källan InfoFinland.fi.
I nödsituationer ringer du nödnumret 112.
När arbetsavtalet gäller tillsvidare har arbetstagaren en fast eller permanent anställning.
För fristående yrkesexamen finns ingen bestämd ansökningstid.
Vad händer i småbarnspedagogiken?
Ibland kan norrsken ses också i södra Finland.
registrerad partner
Enligt Finlands lag ska hinder mot äktenskap prövas om du är finsk medborgare eller permanent bosatt i Finland och uppgifterna om dig finns i befolkningsregistret.
Man kan dock använda bilen tillfälligt innan bilskatten är betald.
I Finland finns många medborgarinstitut (kansalaisopisto) och arbetarinstitut (työväenopisto).
Skolhälsovårdfinska _ svenska
I Helsingfors finns såväl universitet som yrkeshögskolor.
Bouppteckningen ordnas av den person som bäst känner till den avlidnes egendom och skulder.
direkt via lönesystemet om det har en inbyggd teknisk förbindelse till Inkomstregistret eller
Läs mer på InfoFinlands sida Till familjemedlem i Finland.
När perioden har gått kan man ansöka om förlängning för bidraget.
Den förberedande undervisningen varar vanligtvis ett år.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
I vissa enskilda fall kan man avvika från försörjningsförutsättningen om det finns exceptionellt vägande skäl eller om barnets bästa kräver detta.
Hjälp med att få slut på våld
Läs mer om barndagvård, förskoleundervisning och grundläggande utbildning på InfoFinlands sida Utbildning för barn.
Man måste delta i rättegången.
Du måste ansöka om familjeförmåner separat från FPA.
Motion och friluftsliv i Helsingforsfinska _ svenska _ engelska
Sambor kan även upprätta ett skriftligt avtal om hur egendomen ska fördelas om paret går isär.
Om du är medborgare i ett EU-land, Liechtenstein eller Schweiz och vill resa till Finland för en kort period, till exempel på semester, på affärsresa eller för att besöka släktingar, behöver du inget visum.
Läs mer: Tandvård.
I Finland är det vanligt med familjer med en förälder.
02700 Grankulla
Tolkningfinska _ svenska _ engelska
Du kan utnyttja de offentliga hälsovårdstjänsterna i Finland om du har hemkommun (kotikunta) i Finland.
Du kan också leta upp en privat familjedagvårdare som vårdar barnen hemma hos sig, eller anställa en skötare i ditt eget hem.
Du kan också hämta ansökningsblanketten på daghemmet eller vid informationen i stadshuset.
Arbets- och näringsbyråerna i Nylandfinska _ svenska
reparera en enfas skarvsladd (spänning 230 V)
Information om det europeiska sjukvårdskortetfinska _ svenska _ engelska
gymnasiet
Begravningstillstånd
EU-medborgarnas rättigheter som rätten att fritt röra sig och arbeta inom EU:s område och rätten att rösta och ställa upp som kandidat i EU-val
Även kommunerna äger hyresbostäder. De är ofta förmånligare än andra hyresbostäder.
Telefonnumret till den gemensamma telefontjänsten för hälsostationerna i Vanda är 09 839 50 000.
Grundskoleelever får stöd i sitt skolarbete.
Stöd för frivilligt återvändandefinska _ svenska _ engelska _ persiska _ arabiska
Broschyren Makens efternamn och barnets efternamnfinska _ svenska _ engelska
Adjektiven böjs efter dessa genus.
Du kan be om att få tid hos en kvinnlig läkare om du vill.
Besök läkaren före slutet av den fjärde graviditetsmånaden.
I Finland råder religionsfrihet.
Om dina studier i Finland till exempel varar mindre än två år, ska försäkringen täcka sjukvårdskostnader upp till minst 100 000 euro.
Studietiden beror på utbildningsprogrammet och din egen studietakt.
Sysselsättningsutsikter för olika yrken i Finlandfinska _ svenska _ engelska
Det är bra att beakta att parförhållandets form påverkar makarnas rättigheter och skyldigheter, frågor som rör egendom och arv, vårdnad om och underhåll av barn samt adoption.
Den lön som betalas till arbetstagaren är nettolönen (nettopalkka).
Finlands Röda Kors hjälper med att ordna resan till Finland för kvotflyktingens familjemedlemmar när dessa fått uppehållstillstånd.
Du kan diskutera preventivmetoder med skolans hälsovårdare och i vissa kommuner kan skolans hälsovårdare ge dig ett startpaket.
Fråga mer hos FPA.
När du ansöker om en förmån, utreder FPA om du har rätt till FPA:s förmåner.
I vuxenutbildningen avlägger du yrkesexamen som fristående examen.
hittar en arbetsplats eller studieplats,
Du kan också söka till ett separat magisterprogram.
linkkiHälsovårdscentralen:
Du får anvisningar om hur detta påverkar ditt utkomststöd för arbetslösa.
I norra Finland kan temperaturen vara till och med -30 grader.
Mer information om att ansöka om skilsmässa hittar du på justitieministeriets webbplats.
Skolbyrån
För att arbeta måste du ha ett finländskt skattekort.
Du ska ansöka om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut.
Boka tiden via Migrationsverkets elektroniska tidsbokningssystem.
Läs mer om utlänningars rösträtt i Finland på InfoFinlands sida Val i Finland.
I Vanda finns även Finavia Avia College som ger utbildning för olika luftfartsyrken.
Integrationsutbildningen kan omfatta studier i finska, andra studier eller arbetsförsök.
Ansökan om ordningsnummerfinska _ svenska _ engelska
Till exempel FPA och migrationsverket (Maahanmuuttovirasto) beställer i vissa fall en tolk för kunden.
EU-medborgare ska också registrera sig på Migrationsverket.
linkkiEsbo biIdkonstskola:
Om du har problem med alkohol eller andra droger eller spelproblem kan du ta kontakt med A-klinikkaan.
Du kan samtidigt köpa fler andelar i din bostad om du har kommit överens med byggherren om detta.
Preventivrådgivningfinska _ svenska _ engelska
linkkiPyhäjoki kommun:
Reseplanerarefinska _ svenska _ engelska _ ryska
Serviceboendefinska _ svenska _ engelska
Det är möjligt att i enskilda fall avvika från försörjningsförutsättningen, om det finns exceptionellt vägande skäl eller om barnets bästa kräver detta.
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en krismottagning för invandrare.
Boendetiden kan vara från en dag till flera månader.
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Då hyrsvärden väljer hyresgäst får han eller hon enligt lagen inte diskriminera någon exempelvis på grund av etniskt ursprung, religion eller nationalitet.
Besök Migrationsverkets tjänsteställe; du måste styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Alla invandrare har rätt att få grundläggande information om Finland.
Förberedande utbildning för invandrare
Blivande förskolebarn får mer information om detta per post, på dagvårdens webbplats och i lokaltidningen.
Tandvården vid hälsovårdscentralen är avgiftsfri för barn under 18 år.
Läs mer på InfoFinlands sida Våld och Hedersrelaterat våld.
Röda Korset söker försvunna anhöriga och förmedlar meddelanden på krisområden.
Det är inte obligatoriskt att ta studielån.
Därefter kan man fortsätta studierna och avlägga yrkesexamen eller specialyrkesexamen.
I Finland finns också slott som är öppna för allmänheten, till exempel Olofsborg, Åbo slott och Tavastehus slott.
Vanligtvis ansöker man om dagvårdsplats i den egna kommunen.
Deras färdighetsnivå är 1–2.
Naturen i Finland är mångsidig.
Gifta makar av samma kön har rätt att adoptera ett barn och rätt till adoption inom familjen.
Du kan även be om hjälp och råd vid kommunens skuldrådgivning eller socialverk eller en boenderådgivare vid kommunen eller hyreshusbolaget eller till exempel Garantistiftelsen.
Uppehållstillstånd på andra grunderfinska _ svenska _ engelska
Med den här blanketten kan du meddela följande information till myndigheterna:
linkkiEuropeiska unionen:
Svenska språket i Finland.
Var ligger närmaste magistrat, hälsostation eller bibliotek?
Distansgymnasiumfinska
När du flyttar i Finland från en bostad till en annan:
Information om tågtidtabellerna hittar du på VR:s webbplats och på järnvägsstationerna.
När hemvården är regelbunden påverkar dina egna och din makas eller makes inkomster hemvårdsavgiften.
Broschyren Information till asylsökandefinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Läs mer om att bevisa dina språkkunskaper på InfoFinlands sida Officiellt intyg över språkkunskaper.
I Helsingfors finns det flera daghem som drivs av staden och privata daghem.
Motion
Samtalen besvaras av krisarbetare och utbildade frivilliga stödpersoner.
I Finland värdesätts ärlighet.
Fyll i blanketten noggrant och underteckna den.
Då är barnet ca nio månader gammalt.
Om umgänget blir problematiskt
Färdighetsnivåerna i statsförvaltningens språkexaminafinska _ svenska
Rasism och rasistiska brott
Om föräldrarna är gifta kan de välja endera makens efternamn till barnet.
I krissituationer kan du ringa eller åka till jouren.
Ett samboförhållande registreras inte någonstans.
Film om munhälsovårdfinska _ engelska _ somaliska _ arabiska
Läs mer på InfoFinlands sida Rättigheter och skyldigheter för boende.
Tfn (09) 816 45285
till vård av hög kvalitet
Rådgivningen ges av en jurist.
Asylsökande
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
En rörelsenedsättning kan bero på en sjukdom, ett olycksfall eller genetiska orsaker.
Vård utom hemmet betyder att barnet bor någon annanstans än hos sina föräldrar.
Ryska och engelska: 050 325 7173
I ett höghus hittar du ordningsreglerna vanligtvis i trapphuset nära entrédörren.
Om du vistas i Finland utan uppehållstillstånd kan du emellertid bli tvungen att betala för vården.
Vad stadigvarande boende betyder definieras i lagen.
Sambo med en utländsk medborgare
Alla helgons dag firas i början av november.
linkkiKommunbostäder:
Fundera på vilka produktionsmedel eller vilken arbetskraft du behöver.
Mer information om den kommunala ungdomsverksamheten får du hos ungdomsväsendet i din hemkommun.
Ibland finns det i annonsen en utsatt tid då bostaden visas.
Studietillfällena är dock öppna för alla.
Vad är våld?
arbete
När du flyttar ditt stadigvarande boende till Helsingfors, ska du registrera dig som invånare i kommunen.
Ansökan ska lämnas in till FPA senast en månad innan moderskapspenningperiodens utgång och föräldrapenningperiodens början.
Karlebygatan 27, PB 581
Sambor kan ha sådan egendom om vars ägande de inte har en överenskommelse.
linkkiFinansministeriet:
Stadsfullmäktiges sammanträden på Internetfinska
Medborgarinstitutens musikgrupper är öppna för alla.
Bouppteckningshandlingen (perukirja) ska lämnas till skattebyrån senast en månad efter bouppteckningen.
Prövningen tar ungefär en vecka.
Om du söker till ett utbildningsprogram där undervisningsspråket är ett annat än finska eller svenska, beror ansökningssättet på utbildningen.
Boka en tid hos hälsostationens allmänläkare om du till exempel har problem med blödningar eller smärtor i underlivet.
eBiblioteket (eKirjasto) tillhandahåller elektroniska material, såsom böcker, tidskrifter och filmer.
På babyresa - För dig som har fött barnfinska _ svenska _ engelska
Om du har problem eller oklarheter med uppehållstillståndet, kan du ta kontakt med följande instanser för att be om råd:
Du kan bli klient om du flyttat till Finland på grund av familjeband, är flykting, offer för människohandel eller har rätt till en inledande kartläggning.
Vanligtvis är barnets föräldrar dess vårdnadshavare.
Information om skolresestödetfinska _ svenska _ engelska
När du funderar på vilken företagsform du ska välja, är det absolut tillrådligt att du kontaktar företagsrådgivningen.
–15 studeranden och vanligtvis finns det 8–10 undervisningsgrupper.
Fackets ABC-bokfinska _ engelska _ ryska _ estniska
Fråga mer vid din läroanstalt.
Yrkesexamen och specialyrkesexamen ger dig behörighet till ett visst yrke.
Den förberedande utbildningen tar ett läsår och ger beredskap för gymnasiestudier.
som har rösträtt i val till Europaparlamentet och
Information om fackförbundsverksamhetfinska _ svenska _ engelska
I naturhuset Villa Elfvik ordnas utflykter, evenemang och utställningar.
Tfn (09) 5056 357 eller (09) 5056 358
Ateneumfinska _ svenska _ engelska
Broschyren Information om den finska grundskolanengelska _ ryska _ franska _ somaliska _ arabiska
Religiösa seder eller ritualer hör inte hemma på den finländska arbetsplatsen.
Samtidigt får du en ansökningsblankett.
Som bevis duger till exempel ett utdrag ur boenderegistret eller ett hyreskontrakt med bådas namn.
hushållets bruttoinkomster (inkomster före skatt)
Det är bra att ni går till kliniken tillsammans.
Om det behövs kan du få servicerådgivning om användningen av nättjänsterna.
Söndagen är påskdagen och då minns man Jesu uppståndelse.
Ta reda på om du kan skjuta upp andra betalningar för att kunna betala hyran.
Livet kan vara svårt till exempel när man flyttar från ett land till ett annat, har problem på arbetsplatsen, förlorar sin arbetsplats, har problem i familjen, går igenom skilsmässa, förlorar en anhörig, blir sjuk eller när livet förändras på andra sätt.
Mer information hittar du på Helsingfors stads webbplats.
Via tjänsten Religionerna i Finland kan du söka information enligt religionssamfund och ort.
I Helsingfors har papperslösa invandrare rätt att få brådskande och nödvändig vård inom de offentliga hälsovårdstjänsterna.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Borgerliga vigslar förrättas på magistraten.
Du kan få fortbildning eller påbyggnadsutbildning i din egen bransch.
Tfn 045 639 6274 (24h)
Flyttanmälanfinska _ svenska _ engelska
Barnet får utföra lätt arbete några timmar om dagen om det inte skadar hennes hälsa eller skolgång.
linkkiRättsväsendet:
linkkiAnonyma alkoholister, AA:
Yrkesexamen kan även avläggas med läroavtal.
Företagshälsovård
Hur du ansöker om pension till utlandet beror på i vilket land du bor.
Behöver jag ett tillstånd för företaget?
Tjänster av detta slag är bland annat måltidstjänst och transporttjänst.
Du kan delta i yrkesinriktad arbetskraftsutbildning, om
Studerandena inom integrationsutbildningen kommer från tiotals olika länder och undervisningsspråket är finska. En kurs kan ha 8
I dagvården lär barnet känna den finländska kulturen, lär sig det finska språket och verkar i en social grupp.
Längst ner på varje undersida i InfoFinland hittar du en responslänk, via vilken du kan skicka respons som direkt berör innehållet på sidan.
Vård av barnet i hemmet
17 år
Också många arbetsplatser utbildar sina anställda till exempel i användningen av nya apparater eller program.
Om du flyttar ditt stadigvarande boende till Grankulla, ska du registrera dig som invånare i kommunen.
Läroplikten upphör om den inte redan har fullgjorts.
Vasavägen 7
Du måste ansöka om ett nytt uppehållstillstånd på grund av arbete innan ditt uppehållstillstånd för att söka arbete går ut.
Vid Vanda vuxenutbildningsinstitut (Vantaan Aikuisopisto) kan man till exempel skapa konst, handarbeten, laga mat eller dansa.
Om du har en sjukförsäkring i ett annat EU-land, EES-land eller i Schweiz har du rätt till nödvändig sjukvård i Finland.
Vid folkhögskolor kan du även avlägga yrkesexamen.
Rätten till FPA:s förmåner
Böle verksamhetsställe
Fråga bibliotekarienfinska _ svenska _ engelska
Enligt lag har du rätt att välja antingen finska eller svenska som integrationsspråk.
Vissa tv-program kan du titta på avgiftsfritt.
Avdragen beaktas då i din skatteprocent.
Bibliotek
En del arbetsgivare utbildar människor till arbeten hos dem.
Om studeranden har ett annat modersmål än finska eller svenska och saknar tillräckliga språkkunskaper för gymnasiestudierna, kan hen söka till förberedande gymnasieutbildning (LUVA).
Söka tjänster
Merparten av studierna är dock på finska eller på svenska.
linkkiMiljöförvaltningen:
Välkommen!
Utbildning för döva invandrarefinska _ svenska _ engelska
Du kan studera finska som arbetskraftsutbildning.
Den förberedande undervisningen före grundskolan är avsedd för alla de barn med invandrarbakgrund som inte har tillräckliga kunskaper för att klara sig i undervisningen inom den grundläggande utbildningen.
Du själv betalar förmedlingsarvodet endast om du har ingått ett skriftligt uppdragsavtal med bostadsförmedlaren om att söka en bostad åt dig.
På universitet kan man avlägga lägre högskoleexamen på cirka tre år och därefter högre högskoleexamen på cirka två år.
Läs mer: Läkemedel.
