vid tidsbeställningen får du veta hur snabbt du kommer att få vård .
Vanda centrum ligger i Dickursby .
Användarpanelen är öppen för alla som är intresserade av InfoFinland .
du hittar mer information på HRT:s webbplats .
rådgivning för ungafinska
bostadsrättsbostad
vilka hälsotjänster kan du använda ?
på InfoFinlands sida Problematiska situationer i Helsingfors får du information om var i Helsingfors man kan få hjälp med barns och ungas problem , eller vid problem i familjen .
om studeranden har ett annat modersmål än finska eller svenska och saknar tillräckliga språkkunskaper för gymnasiestudierna , kan hen söka till förberedande gymnasieutbildning ( LUVA ) .
senioruniversitetet ( ikäihmisten yliopisto ) är avsett för dem som har fyllt 60 år .
det finska språket och den finländska kulturen och ekonomin utvecklades enormt under Finlands tid som en del av Ryssland .
inga ytterligare begränsningar - Du får inte tillämpa lagliga begränsningar eller teknologiska metoder som juridiskt begränsar andra från att gör något som licensen tillåter .
på mötet kan man komma överens om hur situationen ska lösas .
om du av någon anledning inte till exempel lyckas få en läkartid utanför arbetstiden , ska du komma överens med din chef om att du är borta och hur du ersätter din frånvaro .
en del av tjänsterna i Päihdelinkki finns även på svenska , engelska och ryska .
kvällar och veckoslut är jourmottagningen centraliserad till större vårdenheter .
Rovala @-@ institutets utbildning för invandrare
Lyft fram sådana färdigheter som behövs i uppgiften .
läs mer på InfoFinlands sida Trafiken i Finland .
om du har slutat använda preventivmedel , men en graviditet inte har börjat inom ett år , boka tid på hälsostationen eller hos en privat gynekolog .
en ung som inte är trygg i sitt eget hem kan kontakta Finlands Röda Kors De ungas skyddshus .
som orsak för abort ( abortti ) räcker även att det med tanke på din livssituation skulle vara en alltför stor belastning att föda barnet eller att ta hand om det .
vid mödrarådgivningen ( äitiysneuvola ) följs moderns , fostrets och hela familjens hälsotillstånd under graviditeten .
Adjö .
be om intyget av din arbetsgivare .
om det är svårt eller omöjligt att bo i bostaden under reparationerna , har du rätt att säga upp hyresavtalet eller får nedsatt hyra .
statsförvaltningens språkexaminafinska _ svenska
även våld mot familjemedlemmarna är ett brott .
du kan påvisa dina yrkeskunskaper med ett fristående yrkesprov .
Vanda och hela huvudstadsregionen har goda kollektivtrafikförbindelser .
registreringsintyget över uppehållsrätt för EU @-@ medborgare ( om du är EU @-@ medborgare )
Assistenten kan hjälpa dig till exempel med att laga mat , handla , på din arbetsplats , i dina studier eller dina hobbyer .
om du har din hemkommun i Esbo kan du utnyttja de offentliga hälsovårdstjänsterna .
en myndighet , till exempel en notaries publicus , måste verifiera överenskommelsen .
webbplatsen betjänar även myndigheter i deras Flerspråkiga informationsverksamhet .
företagsverksamheten är din huvudsyssla
våld i hemmet
Anhållan om prövning av hinder mot äktenskapfinska _ svenska _ engelska
då måste samhället ingripa i familjens situation .
du kan även gå till en privat tandläkarmottagning .
vårdbidrag för pensionstagare
information om riksdagsvalfinska _ svenska _ engelska
särskilt lönar det sig att utreda bostadens skick grundligt .
när du väntar barn
dessutom används nationella läroplansgrunder och lokala läroplaner .
om du har en bil måste du teckna en trafikförsäkring ( liikennevakuutus ) .
Finland förlorade båda krigen , men Sovjetunionen ockuperade aldrig Finland .
volontärarbetefinska
linkkiEures @-@ portalen :
dessa ordnas oftast i årskurs nio .
när du söker till ett universitet , får du i allmänhet poäng utifrån studentexamen och inträdesprovet .
hur många år du återbetalar lånet
linkkiFinska ortodoxa kyrkan :
vilka tjänster ditt lands beskickning tillhandahåller beror på lagen i ditt hemland .
Arbetslagstiftningfinska _ svenska _ engelska
meddela alltid
också polisen kan undersöka orsaken till dödsfallet .
integrationsrelaterade socialtjänster
på våren är det mycket svårt att bedöma isens bärkraft och då är det bäst att undvika att färdas på isen .
tidsbeställning på vardagar .
du kan även ringa kristelefonen om du är orolig för en närstående person .
i Esbo finns dessutom familjedagvårdare .
registrering av uppehållsrätt för EU @-@ medborgarefinska _ svenska _ engelska
information om TE @-@ byråns tjänster för invandrare finska _ svenska _ engelska
när föräldrarna skiljer sig ska de komma överens om underhållet av barnet samt om eventuellt underhållsbidrag ( elatusapu ) .
om ditt fostervatten går eller du har tätt återkommande smärtsamma värkar ska du ringa sjukhuset och fråga om det är dags att åka .
om du inte har en bostad eller om du har bostäder på flera kommuners område är din hemkommun den kommun som du själv uppfattar som din hemkommun och som du har någon fast förbindelse till , till exempel genom familjeförhållanden eller arbetsplats .
råd i frågor som rör familjen
jämställdhet mellan män och kvinnor
i vissa fall kan du också få bostadstillägg , till exempel om du studerar på en avgiftsbelagd linje vid en folkhögskola och bor på läroanstaltens internat .
be Fpa om mera information .
det betyder att den som avlägger utbildningen får en arbetsplats hos arbetsgivaren .
Begravningsplatserfinska _ svenska _ engelska
köp hållbara produkter .
du måste betala avgiften samtidigt som du ansöker om fortsatt uppehållstillstånd .
Låt ögonläkaren undersöka dina ögon regelbundet så att eventuella ögonsjukdomar upptäcks i ett tidigt skede .
efter att betänketiden gått ut ska du eller ni ansöka om slutlig äktenskapsskillnad inom ett halvt år .
storleken på hyran varierar beroende på bostadens läge .
på vissa bibliotek ordnas även språkcaféer i det finska språket för invandrare .
tfn 0400.979.175
Friluftsområdenfinska _ svenska _ engelska
7 @-@ 17 @-@ åringar har läroplikt ( oppivelvollisuus ) , d.v.s. skyldighet att avlägga grundskolans ( peruskoulu ) lärokurs .
du kan redogöra för hur du försörjer dig i Finland .
i Helsingfors finns många gymnasieskolor .
Finland är det viktigt att känna till de grundläggande reglerna som gäller i arbetslivet och det finländska samhället .
du kan få hjälp med din rädsla till exempel vid polikliniken för förlossningsrädsla ( synnytyspelkopoliklinikka ) .
Tänk på att arbete som freelancer eller företagare kan påverka din arbetslöshetsförsäkring .
du kan också ansöka om många slags uppehållstillstånd och EU @-@ registrering på internet i tjänsten Enter Finland .
i Esbo finns flera yrkes- och amatörteatrar .
grundläggande utbildning
barnet måste delta i förskoleundervisningen .
information om företagshälsovårdenfinska _ svenska _ engelska
ditt utbildningsbehov
offentliga hälsovårdstjänster tillhandahålls till exempel vid hälsostationer , tandkliniker , rådgivningsbyråer och sjukhus .
arbets- och näringsbyrån väljer studerandena till den yrkesinriktade arbetskraftsutbildningen .
magistraten fattar beslut om registrering av hemkommun .
i Helsingfors beslutas ärenden av stadsfullmäktige .
i början av året skickar staden en anmälan om läroplikt ( oppivelvollisuusilmoitus ) till hemmen .
i Finland fästs stor uppmärksamhet vid arbetssäkerhet .
om du behöver akut tandläkarvård kvällstid eller under veckoslut , kan du kontakta Haartmanska sjukhuset i Helsingfors .
du kan berätta vilka målsättningar du har med jobbsökningen eller vilken specialkompetens du besitter .
på webbplatsen för Suomen lakiopas får du information om vilka handlingar du behöver för bodelningen .
om barnet inte är finsk medborgare måste han / hon ha uppehållstillstånd i Finland .
tfn 075.7575.100
gör videoklippet på något av de språk som används i Infobanken .
Mottagningscentralen betalar mottagningspenning till asylsökande .
vi använder cookies
jourmottagningen tar endast hand om barn med brådskande hjälpbehov .
i Helsingfors finns även ett muslimskt daghem vars verksamhetsspråk är arabiska .
vilka möbler som ingår varierar .
att ansöka om bostadsbidragfinska _ svenska _ engelska
vetenskaplig fortbildning vid universitet
InfoFinland finansieras av staten och samarbetskommunerna .
Familjevård kan även ordnas i den vårdbehövandes eget hem .
flyktingar kan be om hjälp och rådgivning i rättsliga frågor bland annat från Flyktingrådgivningen r.f. eller från rättshjälpsbyråer .
Miessakit rf strävar efter att sörja för mäns välbefinnande och erbjuder sociala aktiviteter och stöd .
databehandling och datakommunikation
Närbiblioteken finns i Björkhagen , Kelviå , Lochteå samt Ullava kyrkby och Rahkonen .
diskriminering på arbetsplatsen
läs mer på InfoFinlands sida Brott .
Seniorernas tjänster , hemvårdfinska _ svenska
om du är under 25 år , kontrollera tilläggsvillkoren för arbetsmarknadsstödet för unga på TE @-@ tjänsternas webbplats .
bokföring
lagar och kollektivavtal reglerar exakt när tidsbundna anställningar får tillämpas .
barnatillsyningsmännen ger även råd till föräldrar som ska skiljas .
i Finland gäller allemansrätten ( jokamiehenoikeus ) .
barns tandvård
fråga om integration på svenska när din inledande kartläggning och integrationsplan görs .
fråga vid socialbyrån om kommuntillägg betalas i din kommun .
vi läser tillsammans i Vandafinska _ svenska _ engelska
om du hemma vårdar en långtidssjuk , handikappad eller äldre familjemedlem kan din hemkommun betala stöd för närståendevård ( omaishoidontuki ) till dig .
Invandrarelever använder i huvudsak grundskolans och gymnasieskolans vanliga tjänster .
du kommer till Finland för att arbeta som tolk , lärare , sakkunnig eller idrottsdomare i högst tre månader utifrån en inbjudan eller ett avtal ;
du kan bo i bostadsrättsbostaden så länge du vill .
Undervisningsgruppen ska ha minst fyra elever .
om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period .
linkkiFinlands flyktinghjälp :
som EU @-@ medborgare kan du ansöka om studieplats vid en läroanstalt som är godkänd i Finland .
det är viktigt att du har tillräckligt med kapital i startskedet .
huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ ryska _ somaliska _ persiska _ arabiska
vaccinationer
i Vanda finns en delegation för mångkulturella frågor ( monikulttuurisuusasiain neuvottelukunta ) som lägger fram propositioner i ärenden som rör invandrare .
Engelsk @-@ finskspråkigt daghemfinska _ engelska
uppehållstillstånd på en ny grundfinska _ svenska _ engelska
bolagsman i ett öppet bolag
om din företagsverksamhet upphör , kan du ansöka om inkomstrelaterad dagpenning ( ansiosidonnainen päiväraha ) vid arbetslöshetskassan .
du kan få arbetslöshetsstöd från och med det datum då du anmälde dig som arbetslös .
linkkiSkatteförvaltningen :
i särskilda fall kan barnet börja skolan senare .
boka tid för vigseln hos magistraten eller tingsrätten i god tid före bröllopsdagen .
du kan ansöka om moderskapspenning om du omfattas av den sociala tryggheten i Finland och varit sjukförsäkrad i Finland , ett annat EU- eller EES @-@ land eller Schweiz oavbrutet i 180 dagar före det beräknade förslossningsdatumet .
Biträdet deltar i asylsamtalet efter sitt eget omdöme .
för registrering av en familjemedlem till en EU @-@ medborgare krävs också att den person som är bosatt i Finland har tillräckliga medel för att försörja sig själv och sin familjemedlem som ska flytta till Finland .
för att du ska kunna få en hemkommun i Finland måste du flytta till och vara stadigvarande bosatt i Finland .
evangelisk @-@ lutherska församlingarfinska _ svenska _ engelska
linkkiStatens rättshjälpsbyrå :
arbete och entreprenörskap
målet är att stödja barnets utveckling och välbefinnande .
hur sorteras avfall ?
om du tänker köpa en bostadsaktie , ta då även reda på vilka renoveringar bostadsaktiebolaget planerar och vad de kostar .
om du vill ansöka om en hyresbostad , fyll i en ansökningsblankett för hyresbostad på Espoon Asunnot Oy:s webbplats .
ni har gemensamma barn eller
utkomststöd kan du få om du inte lyckas få tillräckliga inkomster genom eget arbete , andras omsorg eller på något annat sätt .
du kan ansöka om en delägarbostad med en ansökan riktad till bostadens byggherre .
serviceboende är en boendeform avsedd för sådana personer som behöver kontinuerlig hjälp men inte är i behov av anstaltsvård .
du kan låta utföra ändringsarbeten i ditt hem som underlättar boendet .
Ungdomsgårdarfinska _ svenska _ engelska
med sökmotorn kan du kontrollera var och när du kan avlägga examen .
linkkiUtbildningsstyrelsen :
arbetstagaren kan få ersättning vid ett olycksfall .
mer information får du till exempel på Väestöliittos webbplats eller webbplatsen för kyrkans familjerådgivningscentral .
öppna yrkeshögskolor
på stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang .
du kan även beställa skattekortet via Skatteförvaltningens telefontjänst :
ditt födelseår avgör i vilken ålder du kan få arbetspension .
arbetstiden ska följa arbetslagstiftningen och kollektivavtalet .
adress : Sörnäsgatan 1
penningunderstöd för utländska forskarefinska _ svenska _ engelska
läs mer : högskoleutbildning
när du vill flytta behöver du inte sälja bostaden .
du kan också lämna initiativ och ställa frågor samt kommentera ärenden på finska och på svenska .
motion .
hyresvärden ska meddela hyresgästen om hävandet .
P @-@ EU @-@ tillstånd gäller tills vidare .
legitimation ( till exempel pass )
i Finland råder också yttrandefrihet .
om man redan behärskar de färdigheter som krävs för examen , kan man också avlägga yrkesexamen eller specialyrkesexamen som yrkesprov .
Minimiarbetstiden är vanligtvis 18 timmar i veckan .
Samtalen är konfidentiella .
rätten till en hemkommun i Finland bestäms enligt hemkommunslagen .
val av förlossningssjukhusfinska _ svenska _ engelska
tfn 016.322.8091 eller tfn 016.322.8014
hur ansöker man om en bostadsrättsbostad ?
om du flyttar ditt stadigvarande boende till Esbo , ska du registrera dig som invånare i kommunen .
polisen utfärdar identitetskort .
läs mer : bibliotek
Avsikten är att fadern tar hand om barnet .
föräldrarna kan hjälpa ledarna att utarbeta planen .
om din arbetsgivare är finländare eller om din utländska arbetsgivare har en arbetsplats i Finland , betalar du skatt i Finland .
hyresgästen har rätt att göra detta , om bostadens egentliga hyresvärd godkänner detta .
mer information om motionsrutterna , rastplatser , möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats .
tfn ( 09 ) 839.22133
tjänsten är kostnadsfri .
om du är medborgare i något av de nordiska länderna , ett EU @-@ land , ett EES @-@ land eller i Schweiz och kommer till Finland för att arbeta , behöver du inget uppehållstillstånd .
läs mer : fritid i Esbo
i den finländska kulturen följs dock fortfarande många kristna seder .
1918 inbördeskrig mellan röda och vita
du kan skriva ut blanketten på Migrationsverkets webbplats .
om ett barn blir akut sjukt , ska du ta kontakt med hälsostationen eller jourmottagningen .
statsförvaltningens språkexamen om kunskaper i finska och svenska
allmänt bostadsbidragfinska _ svenska _ engelska
de flesta webbkurser är på finska eller svenska , men det finns även andra alternativ :
om arbetsgivaren säger upp en arbetstagare måste arbetsgivaren ange orsaken till detta .
i Finland finns många föreningar för invandrare .
Helsingfors är Finlands administrativa centrum : där sammanträder Finlands riksdag och där finns ministerierna .
även om Helsingfors växte snabbt , var Esbo ännu länge en fridfull landssocken .
besök läkaren
när du registrerar ditt företag för första gången ska du fylla i en etableringsanmälan och skicka in erforderliga bilagor .
i Esbo finns många olika hotell där man kan bo tillfälligt .
Kompetenscentret Stadin osaamiskeskus ( Stadin osaamiskeskus ) förbereder invandrare för arbetsmarknaden och hjälper dem att hitta ett jobb eller en praktikplats .
du kan söka en jurist till exempel på Finlands Advokatförbunds webbplats , via tjänsten Etsi asianajaja .
använd inte vatten .
det är också viktigt att du bekantar dig med finländare och arbetslivet i Finland redan under studietiden .
avsluta inte samtalet förrän du får lov .
även om du väljer integrationsutbildning på svenska lönar det sig för dig att i något skede även lära dig finska .
begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning .
Kompetenscentret för integration av invandrare stöder arbete som främjar integrationen av invandrare lokalt , regionalt och riksomfattande .
vid tidsbeställningen bedöms vilken slags vård barnet behöver .
du kan till exempel ta vilket som helst namn som du har haft tidigare .
du har rätt att använda arbets- och näringsbyråns tjänster .
du kan även besöka FPA:s kontor .
mer information hittar du på InfoFinlands sida Finska och svenska språket .
Friluftsområdenfinska
brådskande ärenden är till exempel bihåleinflammation , ögoninfektion , ryggvärk , en lindrig urinvägsinfektion , en vaginal infektion eller eksem .
annan orsak
vanligtvis börjar förskoleundervisningen det år då barnet fyller sex år .
barnets officiella adress påverkar också till exempel FPA:s bostadsbidrag .
sambo med en finsk medborgare
svåra livssituationer
du kan få :
om du vill läsa finska eller svenska , läs mer på InfoFinlands sida Finska och svenska språket .
specialyrkesexamina .
om den egna hälsostationen eller det egna sjukhuset inte kan ge patienten vård inom utsatt tid måste de ordna möjlighet för patienten att få vård på ett annat ställe .
flyttanmälan ska alltid göras till magistraten ( maistraatti ) .
om du kommer från ett annat EU @-@ land kan du i vissa fall utnyttja de försäkringsperioder som du har ackumulerat i andra EU @-@ länder .
om du får mer lön än vad du uppgett , överskrids din inkomstgräns .
Arbetsmarknadsstödfinska _ svenska _ engelska
under Stora nordiska kriget år 1710 föll två tredjedelar av Helsingfors befolkning offer till pesten .
Företagsfinland ( via webbplatsen och per telefon )
broschyren jobba i Finland ( pdf , 5,51 MB ) finska _ svenska _ engelska _ ryska _ estniska _ franska _ polska
Biskopsbron 9 B
sambo till en person som fått internationellt skyddfinska _ svenska _ engelska
ett barn eller barnbarn under 21 år som är beroende av din sambo för sin försörjning
vem kan ställa upp som kandidat ?
detta innebär att du på förhand betalar ett penningbelopp som motsvarar några månaders hyra till hyresvärden .
familjerådgivningen betjänar invånarna i Grankulla .
om du vill ansöka om finskt medborgarskap ( kansalaisuus ) kan du påvisa att du har tillräckliga kunskaper i finska eller svenska genom att avlägga den muntliga och skriftliga delen av en allmän språkexamen minst på nivå 3 .
humanistiska och konstnärliga områden
de strävar efter att förbättra dessa minoriteters ställning i samhället .
han eller hon kan således inte hjälpa dig med annat .
Seniorrådgivningenfinska _ svenska _ engelska
den ordnas i daghemmens förskolegrupper .
tjänsten kan också användas av andra invandrare som behöver tillfällig rådgivning i specialfrågor som rör integration .
information om vård av drogproblemfinska _ svenska _ engelska
dessutom ska ditt barn ha en finländsk personbeteckning .
statsborgen kan utgöra högst 20 procent av lånet och högst 50.000 euro .
fråga din arbetsgivare som det ordnas undervisning i det finska språket på din arbetsplats .
Boendeguide för ungafinska
vid arbetarinstitutet kan vem som helst studera .
Återvinningsstationerfinska _ svenska _ engelska
utöver skatt betalar arbetsgivaren försäkringspremier på din lön i händelse av arbetslöshet eller sjukdom .
alla länder har inte en beskickning i Finland .
modern har en finsk personbeteckning .
mer information om att köpa en egen bostad får du på banken eller hos fastighetsförmedlare .
Muslimernas gravkvarterfinska
som studerande betalar du själv vårdkostnaderna om du insjuknar i Finland .
också Helsingfors församlingar har klubbverksamhet .
nyårsdagen 1.1
vid Karleby finska gymnasium anordnas undervisning i finska som andraspråk för invandrare invandrare .
mån kl . 9 @-@ 16 utan tidsbeställning
diskriminering är ett brott .
Sommaruniversitets kurser är avgiftsbelagda för deltagarna .
information om gymnasiestudierfinska _ svenska _ engelska
lämna eller posta blanketten till den dagvårdsenhet där du i första hand söker plats .
äktenskap mellan följande nära släktingar är förbjudet :
observera att utländska handlingar ska vara legaliserade .
Vuxenutbildningsinstitutet ordnar även kurser för invandrare .
gör flyttanmälan senast inom en vecka från din flyttningsdag .
Karleby stads blankett för ansökan om hyresbostad kan fyllas i och skickas in på nätet .
yrkesutbildning efter gymnasiet
studerande
vissa spermiedödande medel kan köpas receptfritt på apotek .
om du till exempel har bokat tid hos en myndighet eller läkaren är det speciellt viktigt att du är på plats i tid .
vanligen består ett hushåll av ett äkta par , sambor eller en familj .
studier i finska språket på Internetfinska _ engelska
hindersprövningen görs på magistraten ( maistraatti ) .
även om du har kommit lagligt till Finland kan din vistelse i landet bli illegal till exempel om du stannar kvar i landet fastän du inte beviljas ett uppehållstillstånd eller om ditt visum eller uppehållstillstånd har gått ut .
till exempel ska lokaler där man säljer livsmedel eller idkar skönhetsvård kontrolleras och tillstånd sökas hos kommunens hälsomyndighet innan lokalerna tas i bruk .
om du till exempel har en krävande hobby eller är sjuk en lång tid kan du avlägga gymnasiet som distansstudier .
barnet kan få minst 20 timmar småbarnspedagogik i veckan eller mer om föräldrarna arbetar eller struderar .
bostadens storlek
Jourmottagningarfinska _ svenska _ engelska
ansökan till yrkesutbildning
skattenummer
linkkiFlyktingrådgivningen r.f. :
linkkiMellersta Österbottens folkhögskola :
ingen får behandlas annorlunda till exempel på grund av kön , ålder , religion eller handikapp .
det finns olika CV @-@ mallar .
här kan du hämta ett skattekort och ett inom byggbranschen obligatoriskt skattenummer .
förlossningen
du kan söka information om rutterna i reseplanerartjänsten ( Reittiopas ) .
den första finskspråkiga ABC @-@ boken ( Aapinen ) ges ut i Finland
under den förberedande undervisningen studerar barnet eller den unga finska och några läroämnen .
att köra bil under alkoholpåverkan är förbjudet enligt lag och det kan ge ett hårt straff .
ersättningen kan vara en ersättning av sjukvårdskostnader och inkomstbortfall i form av dagpenning , olycksfallspension , ersättning för den skada som olyckan har orsakat , rehabilitering eller vid Dödsfall familjepension till de anhöriga .
i Karlebynejden erbjuds olika inkvarteringsalternativ .
åldringar kan använda tjänsterna vid de vanliga hälsostationerna .
i Finland har barn rätt till särskilt skydd och särskild omsorg .
vid problem med din mentala hälsa ska du i första hand kontakta din egen hälsostation eller företagshälsovårdens mottagning .
om ditt land har tillträtt Haagkonventionen ska du begära om ett så kallat Apostille @-@ intyg för din handling .
jag hittar inte en förmånlig hyresbostad .
Uppfostring av barn i Finland ( pdf , 8,08 Mt ) finska _ engelska _ ryska _ somaliska _ kurdiska _ albanska _ burmesiska
Helsingfors evenemangskalenderfinska
när du vill starta ett företag ska du fundera noga på om du har en bra affärsidé .
om du har kommit till Finland som kvotflykting , kan Migrationsverket ersätta kostnaderna för en familjemedlems inresa .
nej : glasföremål , glaskärl , speglar , porslin
telefontjänst : 0295.020.500
anmäla födelsen av ditt barn till myndigheterna i ditt hemland om barnet föds i Finland
läs mer om arbetslöshetskassan på InfoFinlands sida Fackförbund .
linkkiYrkesutövarnas och företagarnas arbetslöshetskassa :
om samborna förvärvar egendom tillsammans ska båda parterna antecknas som köpare och alla kvitton sparas .
Läroavtalsplatsen kan också vara din nuvarande arbetsplats .
om du inte har en sådan handling , kan dina fingeravtryck jämföras med de fingeravtryck som lagrats i uppehållstillståndskortet eller uppehållskortet .
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar .
kom ihåg att företagande även medför risker .
genom att betala en bostadsrättsavgift , som är 15 procent av bostadens anskaffningspris , och därefter varje månad ett rimligt bruksvederlag får man rätt att förvalta över bostaden precis som om den vore en ägarbostad .
företagarkurser
telefonrådgivning : 0295.666.842
arvsskatt
flyktingar kan även kontakta Esbo stads invandrartjänster ( maahanmuuttajapalvelut ) .
företagare i Esbo får även hjälp av Företagarna i Esbo rf .
i Finland finns 40 nationalparker .
när flyktingarna anländer till Finland kommer en anställd från röda Korset till flygplatsen och tar emot dem .
vissa museers samlingar kan du även bekanta dig med på internet .
diskrimineringsombudsmannen kan ge anvisningar , råd och rekommendationer samt hjälpa parterna att åstadkomma förlikning i diskrimineringsfall .
Vailla vakinaista asuntoa ry har ett nattcafé , Kalkkers , som erbjuder bostadslösa en varm plats på natten från höst till vår .
biblioteket producerar även läroböcker för synskadade skolelevers och studerandes behov .
kondomer säljs också till exempel i mataffärer .
Migrationsverket beslutar om du får uppehållstillstånd eller inte .
om du och din granne har en konflikt som ni inte klarar av att själva lösa , kan ni be om hjälp vid grannmedlingscentret Naapuruussovittelun keskus eller hos disponenten .
graviditet kan också förhindras med spermiedödande medel , till exempel p @-@ skum ( emätinvaahto ) eller slidpiller ( emätinpuikko ) , men de är inte särskilt effektiva .
läs mer : studier som hobby
Webbkurs med många hjälpspråksvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
familjeplanering
anvisningar om eftermiddagsverksamhetens klientavgiftfinska _ ryska _ somaliska _ arabiska
på museiförbundets sidor hittar du mer information om dagar med fritt inträde .
sådana hjälpmedel är till exempel datorer och tilläggsutrustning till datorer .
kontrollera ersättningen i ditt kollektivavtal .
linkkiRegionförvaltningsverket :
Ansök om fortsatt uppehållstillstånd elektroniskt i tjänsten Enter Finland eller på Migrationsverkets tjänsteställe .
både myndigheter och vanliga människor deltar i flaggdagarna .
magistraten registrerar dina uppgifter i det finska befolkningsdatasystemet .
barnet behåller sitt tidigare efternamn när föräldrarna skiljer sig .
börjar det år då barnet fyller 7 år
VALMA @-@ utbildningen räcker ungefär ett läsår .
i arbetslivet syns religionens inflytande i de många lediga dagarna som anställda får .
linkkiKarleby kyrkliga samfällighet :
du behöver inte tillstånd av dina föräldrar för receptet .
du betalar avgiften när du lämnar in din tillståndsansökan .
flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum .
information om tandvårdenfinska _ svenska _ engelska
sök tandläkarefinska
Grankulla hälsostation
motiverade skäl för förlängning av visum kan till exempel vara :
kurserna är avgiftsbelagda och de ordnas både dag- och kvällstid .
tolkning för en handikappad är inte det samma som språktolkning .
förmånliga utlandssamtalfinska _ svenska _ engelska
självständiga språkanvändare
ämnen som behandlas på kurserna är till exempel utarbetande av en affärsverksamhetsplan , startande av företagsverksamhet , bokföring , företagsbeskattning , juridiska frågor , marknadsföring , försäljning och kundtjänst .
avgiften är ca 15 procent av bostadens pris .
delta i tävlingen med ditt eget videoklipp !
då är du återflyttare ( paluumuuttaja ) .
information om TE @-@ byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös .
närmare kontaktuppgifter finns på Esbo stads webbplats .
om du på grund av skada eller sjukdom inte kan arbeta kan du få invalidpension ( työkyvyttömyyseläke ) .
den finansieras med skattemedel och är därför förmånligare för familjerna .
när äktenskapets lagliga villkor uppfylls kan ett par gifta sig .
när du går till magistraten ska du ta med dig
i Finland äter man lunch tidigare än i många andra länder .
linkkiTjänstemannacentralorganisationen STTK :
linkkiFinland @-@ samfundet :
därefter övergår eleven till en vanlig klass .
på många metrostationer kan du parkera din bil gratis för att fortsätta resan med kollektivtrafiken .
Finland som en del av Sverige och Ryssland
mer information om anmälan får du på Utbildningsstyrelsens ( Opetushallitus ) webbplats .
att ansöka om partiell sjukdagpenningfinska _ svenska _ engelska
körkort
utlänningar som bor stadigvarande i Finland och som har fyllt 18 år har rätt att rösta i kommunalval .
tidsbokning och rådgivningfinska _ svenska _ engelska
Karlebystödfinska _ svenska
ofta ingår rättsskyddsförsäkringen i hemförsäkringen .
på motionsslingorna kan man springa på somrarna och åka skidor på vintrarna .
du kan söka till dessa utbildningar i den kontinuerliga ansökan året om eller i den gemensamma ansökan till andra stadiet .
vid behov kan du försöka förhandla om att avsluta hyresavtalet tidigare .
betalningen av utkomststöd påverkas av alla dina inkomster och tillgångar .
Mödrahemmets tjänster är avsedda för personer som har hemkommun i Finland .
nattetid kl . 22 @-@ 8
Badhuset / simhallen Vesihiisi
Munhälsovårdenfinska _ svenska
läs mer om Inkomstregistret och om att anmäla löner på Inkomstregistrets webbplats .
vid hälsopunkten Daalia ges vägledning och rådgivning för personer över 65 år om diet , motion och livsstil .
Studiebostäderfinska _ engelska
information om Finlands historiaengelska _ ryska _ franska _ spanska _ tyska _ portugisiska
identitetsbevis ( till exempel pass )
du får studiehandboken till exempel på bibliotek eller Vandainfo samt i elektroniskt format på Vanda stads webbplats .
det grundläggande utkomststödet täcker även utgifter för hobby- och rekreationsverksamhet , avgifterna för barndagvård och för skolbarns morgon- och eftermiddagsverksamhet samt nödvändiga kostnader för flytt .
arbetsgivaren har skyldighet att :
du ska söka med en separat ansökan t.ex .
uppsägningstid
en del privata läkarstationer erbjuder denna tjänst . ett hembesök av en privatläkare är dock dyrt .
Jämför olika mäklarbyråers priser på förhand .
mer information om den förberedande undervisningen för invandrare får du av stadens undervisningstjänster .
Yles radiokanal Mondo erbjuder radioprogram på engelska och många andra språk .
uppehållstillstånd för studerande beviljas högst för två år i taget .
Gränskontrollmyndigheten eller polisen registrerar dig som asylsökande , antecknar uppgifter om dig och tar dina fingeravtryck .
flerfaldigt medborgarskap
man kan resa nästan över allt i Finland med tåg eller buss .
barns och ungas problem
studieplats
är jag offer för människohandel ?
föreningen för bostadslösafinska _ engelska
faderskapet kan erkänns redan under graviditeten vid mödrarådgivningsbyrån eller efter barnets födelse hos barnatillsyningsmannen i den egna kommunen .
läs mer : hälsovårdstjänster i Finland .
flyktingar och asylsökande samt andra utlänningar kan söka hjälp och råd i frågor kring uppehållstillståndet hos Flyktingrådgivningen rf .
när du söker asyl utreder Migrationsverket samtidigt om du kan få uppehållstillstånd på någon annan grund .
Idrottstjänsterfinska _ svenska _ engelska
kontrollera regelbundet att vattenledningarna i ditt hem inte läcker och att det inte rinner ut vatten från hushållsapparaterna på golvet .
du kan hämta en personbeteckning och samtidigt registrera ditt tillfälliga boende i den närmaste magistraten ( maistraatti ) eller skattebyrån ( verotoimisto ) .
då du kommer till sjukhuset ska du använda centralsjukhusets huvudingång kl . 7 @-@ 20 och övriga tider bör du använda den gemensamma jourens / poliklinikens dörr .
mer information får du via tjänsten Helsingforsregionen.fi .
förskoleundervisningen börjar i augusti och ansökningstiden är i januari .
bostäder för bostadslösafinska
information om skyddshem och mödrahemfinska
om du inte får hjälp av din förman ska du ta kontakt med arbetsplatsens arbetarskyddsfullmäktige ( työsuojeluvaltuutettuu ) eller förtroendeman ( luottamusmies ) .
det är inte tillrådligt att säga upp hemförsäkringen under tiden då du bor i bostaden .
när man talar om lön avser man oftast bruttolönen ( bruttopalkka ) från vilken skatter och personalbikostnader dras av .
de annonseras inte ut öppet , utan arbetsgivarna söker arbetstagare via sina egna nätverk .
parförhållandet registreras på magistraten .
du hittar information om arbetstagarens rättigheter och skyldigheter i Finland på InfoFinlands sida arbetstagarens rättigheter och skyldigheter .
dessutom erbjuder även privata musikskolor och -institut undervisning .
vissa inträdesprov omfattar förhandsuppgifter .
Skattefinska _ svenska _ engelska
om du har hemkommun i Finland.har du rätt att få dessa undersökningar gjorda .
du kan ansöka om stöd för närståendevård hos socialbyrån i din hemkommun .
om du misstänker att barnets hälsa eller säkerhet äventyras när barnet träffar den andra föräldern ska du meddela detta till socialmyndigheter .
finska 029.497.000
observera att tull- och skattefriheten för flyttsaker inte gäller alkohol eller tobaksprodukter .
mer information om jämställdhet hittar du på InfoFinlands sida Jämställdhet och likabehandling .
tandvårdens jourmottagning kvällar och veckoslutfinska _ svenska _ engelska
är du studerande lönar det sig att ansöka om en studentbostad då dessa vanligen är förmånligare än andra hyresbostäder .
Mannerheims barnskyddsförbund MLL
om du planerar adoption inom familjen ska du kontakta socialbyrån i din hemkommun .
om förlossningen kan utgöra en risk för din hälsa
rådgivning för att motarbeta diskriminering
området hade en direkt förbindelse till Helsingfors .
stadslotsen har jour i områdets bibliotek vissa veckodagar och klockslag .
fyll ansökan i tjänsten Studieinfo.fi .
bostäder säljs av privatpersoner , fastighetsförmedlingar och byggherrar .
på Väestöliittos webbplats hittar du information om olika preventivmedel .
läroanstalten kan kontrollera att du har tillräckliga språkkunskaper för studierna .
Basfakta
det betjänar invandrare som är bosatta i Rovaniemi och annorstädes i Lappland .
du hittar urvalet av språk i tjänsten i menyn uppe på sidan .
du kan lämna in ansökan om skilsmässa till tingsrätten i din egen eller din makas / makes hemkommun .
läs mer :
Rehabiliteringspenningfinska _ svenska _ engelska
möbler och andra husgeråd
hur ansöker jag ?
lån som beviljas av banker eller Finnvera är vanliga finansieringskällor för många nya företagare .
du ska besöka tjänstestället inom tre månader efter att ha gjort ansökan .
- Om du vill kan du även lista dina publikationer eller arbetsprov .
dessutom ska du ha hemkommun i Finland den 51:a dagen före valdagen .
om du inte är medborgare i något av Europeiska unionens medlemsländer , ett EES @-@ land eller i Schweiz och vill driva ett företag i Finland , behöver du ett uppehållstillstånd för företagare .
om du ska utföra säsongsarbete i Finland behöver du ett säsongsarbetstillstånd .
Mellersta Österbottens och Österbottens rättshjälpsbyrå
läs mer : barn vid skilsmässa
du får mer information om att legalisera officiella handlingar vid magistraten eller beskickningen för ditt eget land i Finland .
senare kan du köpa hela bostaden så att den blir helt och hållet din egen .
vem kan få en bostadsrättsbostad ?
information för utvecklingsstörda och anhörigafinska
största delen av verksamheten på ungdomsgårdarna är gratis .
det är avgiftsfritt .
om du har en hemförsäkring , och din bostad blir skadad till exempel vid en brand eller till följd av en vattenskada , kontakta då genast ditt försäkringsbolag .
vi har samlat kontaktuppgifter till myndigheterna på InfoFinlands sida Ring och fråga om råd .
om du ämnar flytta utomlands från Finland för två år , till exempel på grund av arbete eller studier , kan du ansöka hos Migrationsverket om att ditt uppehållstillstånd inte återkallas .
detta måste du emellertid alltid komma överens om med hyresvärden .
linkkiMellersta Österbottens sommaruniversitet :
religionsfrihet och religionsutövande i Finland
efter grundskolan ( peruskoulu ) , d.v.s. efter grundstadiet fortsätter studerandena till läroanstalter på andra stadiet ( toisen asteen oppilaitos ) .
tfn ( 09 ) 8789.1344
