��      ]�(�numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����i4�����R�(K�<�NNNJ����J����K t�b�C<      �      �  :   M     (      x   "   �        �t�bhhK ��h��R�(KK��h�CD1        A   �     K  ?      
   &           F         �t�bhhK ��h��R�(KK��h�C4      J   a      �  &                    �t�bhhK ��h��R�(KK��h�C8   �         L  �      �   ]   )   d   �         �t�bhhK ��h��R�(KK��h�C8�     N  �     8   E  y      �               �t�bhhK ��h��R�(KK��h�C4#   !      x   (      :   %        �        �t�bhhK ��h��R�(KK��h�CT   b      �   G   �        J   �   <     �         .                  �t�bhhK ��h��R�(KK��h�CP   (   -   x               �     [      8   �      �     o         �t�bhhK ��h��R�(KK��h�CL      5   �   9   �   �  &      U     �   
   �  *     �        �t�bhhK ��h��R�(KK��h�C4   .   �           �  �  =     @         �t�bhhK ��h��R�(KK��h�C�  �   �  �
        �t�bhhK ��h��R�(KK��h�C0�  �
     �  �     
      :   O        �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�CD      =         =  M  *         
  8   �  :   O        �t�bhhK ��h��R�(KK	��h�C$      )   F  >  
   &        �t�bhhK ��h��R�(KK��h�C<      '     �  
   ?           
   A   }         �t�bhhK ��h��R�(KK��h�C`	  (  �     p            �             �     $   �     @     $  	        �t�bhhK ��h��R�(KK&��h�C�      )   \  N  "         �        
         O  �  j   �  �       �      �           �   �     �  �      �              �t�bhhK ��h��R�(KK��h�CdA        �
  �
                   �         �
     �              �  F        �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C    >   
  L   "   �        �t�bhhK ��h��R�(KK��h�CX�
     �
                 �   �  �   "   @      X      e                �t�bhhK ��h��R�(KK��h�C�     X      �t�bhhK ��h��R�(KK��h�CD      ~      P     �     �
  @   '      "   Q  �        �t�bhhK ��h��R�(KK��h�C4M     
   R  y         �   �              �t�bhhK ��h��R�(KK��h�C<�      �  �     �
     �     0   <   "   �
        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD      2        �  �   �   "   �       '  O  7         �t�bhhK ��h��R�(KK��h�C P  5   �   3  :   +          �t�bhhK ��h��R�(KK��h�C0      &   �   �            G  ]  �     �t�bhhK ��h��R�(KK��h�C              �t�bhhK ��h��R�(KK
��h�C(�  �       B       �        �t�bhhK ��h��R�(KK��h�C   �  �  �         �t�bhhK ��h��R�(KK��h�C/   "   �      �t�bhhK ��h��R�(KK��h�C�      �t�bhhK ��h��R�(KK��h�C4   �  �  $     �     l   9     7         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK	��h�C$H   �     (  S  -   �        �t�bhhK ��h��R�(KK	��h�C$)     �   *   Q     �        �t�bhhK ��h��R�(KK��h�C0   X   �   )   H      V   C    m        �t�bhhK ��h��R�(KK��h�CD        �          �t�bhhK ��h��R�(KK��h�CP  j      	         �t�bhhK ��h��R�(KK��h�C�   E  	         �t�bhhK ��h��R�(KK	��h�C$T        �                 �t�bhhK ��h��R�(KK��h�C4U  4     A   F     *     �
  +   n         �t�bhhK ��h��R�(KK��h�C<"   �              (      <      �     G        �t�bhhK ��h��R�(KK��h�C\$     �     +         5      V        �      �   :            O           �t�bhhK ��h��R�(KK��h�C�   �     �      �     �t�bhhK ��h��R�(KK��h�C�  �  	      	         �t�bhhK ��h��R�(KK	��h�C$�     L  �      �  �         �t�bhhK ��h��R�(KK��h�CH      O         Y      Q      Q     Q      x              �t�bhhK ��h��R�(KK��h�C`      0   R  <   "      �
  )   
               )               G     )        �t�bhhK ��h��R�(KK��h�C W     �
  	      	         �t�bhhK ��h��R�(KK��h�C\
   �     �     F   '      H     %        *  �      *         �   �         �t�bhhK ��h��R�(KK��h�C@)     /      �   L   G   �     0      �     �        �t�bhhK ��h��R�(KK��h�CI           �t�bhhK ��h��R�(KK��h�C8#   !      �     �  ?      
   3   6            �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK%��h�C�X  �        �  a  �      �     �  
   Z                    
   �        M   �      �
              �  >     �         �t�bhhK ��h��R�(KK��h�CT"           /      �   z   �     "     �
     /      ^  z           �t�bhhK ��h��R�(KK	��h�C$+  �   �  �
  �      �         �t�bhhK ��h��R�(KK��h�C�  Y  �      Z       �t�bhhK ��h��R�(KK��h�C          H   o            �t�bhhK ��h��R�(KK��h�C�  �
  [     �t�bhhK ��h��R�(KK��h�C0#   !         (      
   3   6   �        �t�bhhK ��h��R�(KK��h�C      �  �        �t�bhhK ��h��R�(KK��h�Cb     �      �        �t�bhhK ��h��R�(KK��h�C       �                  �t�bhhK ��h��R�(KK��h�Cd      ~      ,     �
  &      �   -   �   �     �    �                          �t�bhhK ��h��R�(KK
��h�C(      &   \     �  
   c        �t�bhhK ��h��R�(KK��h�C            �t�bhhK ��h��R�(KK��h�C8d  S  \   �  ]     �      �  �  �           �t�bhhK ��h��R�(KK��h�C�  	         �t�bhhK ��h��R�(KK��h�C<�  (   %      R  H        �                    �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0   '      .   
   e     5     y        �t�bhhK ��h��R�(KK��h�C{         S   4      �t�bhhK ��h��R�(KK��h�C~   +           �t�bhhK ��h��R�(KK	��h�C$      f     �      �  f     �t�bhhK ��h��R�(KK��h�C@  &   N   ^         /      �     J     &        �t�bhhK ��h��R�(KK��h�C0�  �     T  
   �     �     @         �t�bhhK ��h��R�(KK��h�C\�   f     g  (  �   )   _     /      �      �                   �
        �t�bhhK ��h��R�(KK��h�CL   �    
   \   H   �        �     \   H   _  %      �        �t�bhhK ��h��R�(KK
��h�C(-   K     ;      �     �        �t�bhhK ��h��R�(KK��h�C0�     �        �
  M     �   �
        �t�bhhK ��h��R�(KK��h�C0      -   �   '     6  
   �            �t�bhhK ��h��R�(KK��h�C   &   N      �      �t�bhhK ��h��R�(KK��h�CH      5   !      �           �   �         �               �t�bhhK ��h��R�(KK��h�C@   
   �   �   -  �   :              �  q   �        �t�bhhK ��h��R�(KK	��h�C$�     z      ,         �      �t�bhhK ��h��R�(KK��h�C<         �      �     �
     �     �  
   �     �t�bhhK ��h��R�(KK��h�C`     �     �         �t�bhhK ��h��R�(KK��h�C,     �t�bhhK ��h��R�(KK��h�C@U   t   
   $   �     �
     U       S     +         �t�bhhK ��h��R�(KK��h�CDV     �     .    �     >   �  *                     �t�bhhK ��h��R�(KK��h�C �   [      �     �          �t�bhhK ��h��R�(KK
��h�C(   �  �      �        �        �t�bhhK ��h��R�(KK��h�C<      z     a     L  z  {  a       b        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK	��h�C$�  h  H   R      �           �t�bhhK ��h��R�(KK��h�CD�   7  (   2      
  �  �   s  :   ?  �  Q     �        �t�bhhK ��h��R�(KK��h�C8"   m   G   �      -  �   �  /  i              �t�bhhK ��h��R�(KK��h�CT   (   <      �  
   �      (        �  �          |      �         �t�bhhK ��h��R�(KK��h�C 2     �
  	      	         �t�bhhK ��h��R�(KK��h�CTj     �  �        �  M  �   �      �
       �   �  }      �
        �t�bhhK ��h��R�(KK��h�CH      w   �       �   �             &  *      �        �t�bhhK ��h��R�(KK��h�C4N  c   I  
   �  F      �                �t�bhhK ��h��R�(KK��h�C`        �     �t�bhhK ��h��R�(KK��h�C0�     �     =         �  G   P        �t�bhhK ��h��R�(KK��h�CO              �t�bhhK ��h��R�(KK��h�Cx   �  9     �  g  �   �  (      !      \         �     �     c  
      k  �     �
  �
           �t�bhhK ��h��R�(KK��h�C �   "   T     �      �     �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK#��h�C�   5   �           8   �                    �      �  P  
   c                 �   �     �
     �             �t�bhhK ��h��R�(KK	��h�C$1   #       *      �  /         �t�bhhK ��h��R�(KK��h�C          �              �t�bhhK ��h��R�(KK��h�CD            �  G      �        =      [   G   H        �t�bhhK ��h��R�(KK��h�CP   %   0  �     2   z  W        �     1        %   �  �        �t�bhhK ��h��R�(KK��h�C �      f   �             �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C!      �        �t�bhhK ��h��R�(KK��h�C         .   �        �t�bhhK ��h��R�(KK��h�C  E      �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C@   (   #   !      X     k   
   3   6   2              �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C/      8     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C �  )                   �t�bhhK ��h��R�(KK��h�CT�  �     N   �      �  �  �     J  
   C   �  -   �                �t�bhhK ��h��R�(KK��h�C     �     �     �t�bhhK ��h��R�(KK��h�C   �     `   �     �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK	��h�C$
     �  %     Q          �t�bhhK ��h��R�(KK��h�C`      R  �
       �   R         �  9   �  �        :            �  �        �t�bhhK ��h��R�(KK��h�CL   X   '   -   H   A   F     L  %   .           �     �        �t�bhhK ��h��R�(KK��h�CP2                �   �         .      S     �        �        �t�bhhK ��h��R�(KK��h�C@�                   �   �        �              �t�bhhK ��h��R�(KK��h�C          W        @      �t�bhhK ��h��R�(KK��h�C%      ~               �t�bhhK ��h��R�(KK��h�C`   l               l      A           �
     0   <      d     %   �          �t�bhhK ��h��R�(KK��h�CD�  �     q   .    V   2      e  C   h   H   B   3        �t�bhhK ��h��R�(KK��h�C  	      	   K      �t�bhhK ��h��R�(KK��h�C4K       �       �      �     9        �t�bhhK ��h��R�(KK
��h�C(!      	        	      	         �t�bhhK ��h��R�(KK��h�C �
        	      	         �t�bhhK ��h��R�(KK��h�C`4                �   �         0   �  �  -                        .         �t�bhhK ��h��R�(KK��h�Clf  
     �  	      	      	   K   	   �   	   �   	     	   I  	   �  	   U  	   �  	   �      �t�bhhK ��h��R�(KK��h�C0      �  �
     �   >        �         �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6            �t�bhhK ��h��R�(KK��h�C0
   �   F   '   !           �  �         �t�bhhK ��h��R�(KK
��h�C(�      /         	      	         �t�bhhK ��h��R�(KK��h�C!            �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C<        {      �     )  +      |      �         �t�bhhK ��h��R�(KK��h�CP   (   �  3  "   @        T     8   �     �  �                 �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�CLY  h     �     h        O     g              �  U        �t�bhhK ��h��R�(KK��h�C�      �   0   <   r      �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�CL         9   9  7      5   �     M   �      �  "   $           �t�bhhK ��h��R�(KK��h�C8   (   �     *      �  +        G   t         �t�bhhK ��h��R�(KK��h�C�
     	      	         �t�bhhK ��h��R�(KK$��h�C�            �  4      �     �               Z        0      k            �
           $        �   �               �t�bhhK ��h��R�(KK��h�C8      �  h     
   �  (   %   )   �           �t�bhhK ��h��R�(KK	��h�C$   [  :     ?  �
  �        �t�bhhK ��h��R�(KK��h�CT   �
     J    /   &   %   �   5     �  |  
   �        "   �         �t�bhhK ��h��R�(KK	��h�C$H   �        �   �           �t�bhhK ��h��R�(KK ��h�C�            i  
   4  P  �   +      �  �     C      6     P               \  L   y      ]  �         �t�bhhK ��h��R�(KK	��h�C$   �      L                 �t�bhhK ��h��R�(KK��h�C@   �   �
  '   �        V         i  �             �t�bhhK ��h��R�(KK��h�C,   f   �    )   �   �      �
        �t�bhhK ��h��R�(KK��h�Cl:   ?  �  Q     �  (      M      +            j  �     �   �
     �  A  �   k  �
        �t�bhhK ��h��R�(KK��h�C<      �        �   j   �     �   9     7         �t�bhhK ��h��R�(KK��h�C    	      	         �t�bhhK ��h��R�(KK��h�C@  �  c                          f   A   �
        �t�bhhK ��h��R�(KK��h�CH           &  *      �        �       �   �  w         �t�bhhK ��h��R�(KK��h�C0�  �  �     �  �        �           �t�bhhK ��h��R�(KK��h�C�     �  r      �t�bhhK ��h��R�(KK��h�CD      �  5   <               �  &      �   j  /        �t�bhhK ��h��R�(KK
��h�C(�   q   7     �     `  �
        �t�bhhK ��h��R�(KK��h�C,      �      P     �   
           �t�bhhK ��h��R�(KK��h�C   	         �t�bhhK ��h��R�(KK��h�C@"   �   �   2        G   %  K  D      �   l          �t�bhhK ��h��R�(KK��h�C �           V     u      �t�bhhK ��h��R�(KK��h�CD�  a     �   W  �     �   f   W  >      w   =            �t�bhhK ��h��R�(KK��h�CX            N  �                             5      �  �  �        �t�bhhK ��h��R�(KK
��h�C(      �           J  E         �t�bhhK ��h��R�(KK��h�C!          �t�bhhK ��h��R�(KK��h�CX      0   �      8   �  �  �  �
     �     "     V     �      �         �t�bhhK ��h��R�(KK!��h�C�   �   �     0   4   -      �      �      �         t        6        l           y   �  �   W              �t�bhhK ��h��R�(KK��h�Cp      M     �t�bhhK ��h��R�(KK��h�C�   �           �t�bhhK ��h��R�(KK��h�Cb     �t�bhhK ��h��R�(KK��h�CL   �    �     7   �
     �     g      �     �     �        �t�bhhK ��h��R�(KK��h�C8#   !      �                               �t�bhhK ��h��R�(KK��h�C1   #       �         �t�bhhK ��h��R�(KK��h�C@1   #         }     o   
   3   6   7  }     o         �t�bhhK ��h��R�(KK	��h�C$�
           C   
   �        �t�bhhK ��h��R�(KK
��h�C(   m  )  �   *   Q     �        �t�bhhK ��h��R�(KK��h�C4      �  �     �      �                 �t�bhhK ��h��R�(KK��h�C  X     �t�bhhK ��h��R�(KK��h�C<�         e  +   
   �     �      v      �         �t�bhhK ��h��R�(KK��h�C �         �  �           �t�bhhK ��h��R�(KK��h�C<      -   �   8        �   o      �      n        �t�bhhK ��h��R�(KK��h�CY            �t�bhhK ��h��R�(KK��h�C4      �
  8  �
     Z       �  �        �t�bhhK ��h��R�(KK��h�CT*      �           �              )        n        ,           �t�bhhK ��h��R�(KK��h�Co     �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6   �        �         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C0�  �  �   �  �       [     �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�Cp^   \        a   �      d   ]     0   !      d   �     ^        �   p     �                  �t�bhhK ��h��R�(KK��h�C0      n      \  L   y                  �t�bhhK ��h��R�(KK	��h�C$�      )   v         0        �t�bhhK ��h��R�(KK��h�C0D   (   �  o  �   "   �     �   �          �t�bhhK ��h��R�(KK��h�CT   ]   �   &      =         �   ~     �  $        t      �           �t�bhhK ��h��R�(KK��h�C8#   !      �  ?      
   3   6   �             �t�bhhK ��h��R�(KK	��h�C$           �
              �t�bhhK ��h��R�(KK��h�C|   L     `     �  �       7   m  �
  7      �
          `     �       9  7      �  �  �        �t�bhhK ��h��R�(KK
��h�C(B    #             +         �t�bhhK ��h��R�(KK��h�C\   <      �           P        �     ,      @      X      e              �t�bhhK ��h��R�(KK��h�C8   ]   �   >      �           �
     H        �t�bhhK ��h��R�(KK��h�CT   S   G         
           $  �  '   �     *           �
        �t�bhhK ��h��R�(KK��h�C�  O      �t�bhhK ��h��R�(KK��h�CHq           %  +         S      q              @         �t�bhhK ��h��R�(KK��h�C 1   #       �     _        �t�bhhK ��h��R�(KK
��h�C(   �  k    
   ,               �t�bhhK ��h��R�(KK��h�C<p     �  �   �  �  �      �  "   �   �   �        �t�bhhK ��h��R�(KK��h�C    @   '   �             �t�bhhK ��h��R�(KK��h�C,   "   �   n        	      	         �t�bhhK ��h��R�(KK��h�C@
   &     �      �  �  +        c   �     �
        �t�bhhK ��h��R�(KK��h�C,      �      �  �  �  �   �
        �t�bhhK ��h��R�(KK��h�CL`  �  :              d   �  ^     �     D   �  N  7         �t�bhhK ��h��R�(KK��h�CP   ?   1     #   !      E      4      �  
   �     q  q   _        �t�bhhK ��h��R�(KK��h�C<                  �     9   '     $   E         �t�bhhK ��h��R�(KK��h�CP   .   r  C      �   O     �     �     u     :  �              �t�bhhK ��h��R�(KK	��h�C$(  s  (   J     I           �t�bhhK ��h��R�(KK��h�CT
   3   6   )  ?   �   �   r   '   !      \         �     �               �t�bhhK ��h��R�(KK��h�C,�         0   [      �              �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6   �     �  m         �t�bhhK ��h��R�(KK��h�CXR  M        �     ]     �   �                 ,            �        �t�bhhK ��h��R�(KK
��h�C(               a  j   �
        �t�bhhK ��h��R�(KK��h�CD#   !      �  �  ?      
   3   6              �        �t�bhhK ��h��R�(KK��h�C�         �     u      �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   �  "   �         �t�bhhK ��h��R�(KK��h�CL�   �
     �   �              !  �      "     �      #        �t�bhhK ��h��R�(KK��h�CT         2                      +      ;  +         o  <        �t�bhhK ��h��R�(KK��h�C8         �         P   +  ^   =  b  *        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C 1   #       `     t        �t�bhhK ��h��R�(KK��h�C<u  �
     $         %  &  �        '  (        �t�bhhK ��h��R�(KK��h�C,   (   T   )     �        v        �t�bhhK ��h��R�(KK
��h�C(      *  +  +         ,        �t�bhhK ��h��R�(KK��h�Ct�        �             %   w  �      �  �         �  �   �  C  !  >     8        -        �t�bhhK ��h��R�(KK��h�C<�
     x       c  	   U  	   �   	   �  	         �t�bhhK ��h��R�(KK��h�C+     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CL
   3   6   �
     �
        '   !      �        �              �t�bhhK ��h��R�(KK��h�C<
   �        e  �
  �
  �   �      ?             �t�bhhK ��h��R�(KK��h�C0�     �     d  <            .        �t�bhhK ��h��R�(KK	��h�C$%      �     �  �           �t�bhhK ��h��R�(KK
��h�C(   �  �   �          �           �t�bhhK ��h��R�(KK��h�C/  	         �t�bhhK ��h��R�(KK��h�Ce     �     �t�bhhK ��h��R�(KK��h�C4*           '   �  H   �     8   S        �t�bhhK ��h��R�(KK��h�CT      �      �  C         �   +     "  g            �              �t�bhhK ��h��R�(KK
��h�C(
   �  6   '   !         ,        �t�bhhK ��h��R�(KK��h�CD   @         �  �  G   k              W              �t�bhhK ��h��R�(KK��h�C0]   P     %         ;      �   �        �t�bhhK ��h��R�(KK��h�Cb   #   "   $            �t�bhhK ��h��R�(KK
��h�C(      -      :  g   0  p        �t�bhhK ��h��R�(KK��h�C4'   !      \         �     �               �t�bhhK ��h��R�(KK��h�C a        	      	         �t�bhhK ��h��R�(KK��h�C4   $   k      X         �   Q  �   �        �t�bhhK ��h��R�(KK��h�C      y  �   �      �     �t�bhhK ��h��R�(KK��h�C4      ,  "   T     :     $   �  �        �t�bhhK ��h��R�(KK
��h�C(I     :   `   3  �      �         �t�bhhK ��h��R�(KK��h�C0�   _        f  �   
   A  �  z        �t�bhhK ��h��R�(KK��h�C g  �  �
        �         �t�bhhK ��h��R�(KK��h�C0�  �     �                 ^        �t�bhhK ��h��R�(KK��h�C</            S   X  i   ,            0   0        �t�bhhK ��h��R�(KK
��h�C(X   �   p  9   W  7     �        �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C �     �  	      	         �t�bhhK ��h��R�(KK��h�C�   -     �t�bhhK ��h��R�(KK��h�C1  	      	         �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�C
   ,   �
  2   �        �t�bhhK ��h��R�(KK��h�C<      �        {  �        �   2     "        �t�bhhK ��h��R�(KK��h�C<H        h     u            3  C   
            �t�bhhK ��h��R�(KK��h�CP      ~         +  &      �   �     �  �   $   .  n      L         �t�bhhK ��h��R�(KK��h�CD   /            |  �      q          �     �        �t�bhhK ��h��R�(KK��h�C1   #       i        �t�bhhK ��h��R�(KK
��h�C(      �      �
  @  N  �         �t�bhhK ��h��R�(KK	��h�C$�   �   �  A  :        �     �t�bhhK ��h��R�(KK��h�Cl   2   J     :  �     �   �  B     >   2   �   �  C   �   7      A  :   �   �     �         �t�bhhK ��h��R�(KK
��h�C(�   >   4  c   
   _      �         �t�bhhK ��h��R�(KK��h�C!         	         �t�bhhK ��h��R�(KK��h�CX%   �          j     �        k     R                    /         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CD4  �     \   �  �      �   +      �      -  d   �        �t�bhhK ��h��R�(KK��h�C5  	      	         �t�bhhK ��h��R�(KK#��h�C�         �   G      t  &      =      n     �     Y      O   
   _      �     �   �        
   �     �     �        �t�bhhK ��h��R�(KK��h�C�
     �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�CL
   t   C  2            "     F     k      l        +         �t�bhhK ��h��R�(KK��h�Ch      ;      �   �      �  R            
  0  4      �        +  4      m           �t�bhhK ��h��R�(KK	��h�C$      }           �        �t�bhhK ��h��R�(KK��h�C`   r     �  +     �  �     �  L         2         �       �
     e        �t�bhhK ��h��R�(KK��h�CL
        �
  6  n     �     �
  �     �     ?      !         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C4D      )   2     �  �      �     �        �t�bhhK ��h��R�(KK��h�C@m     Y      �     )      
   �   �     +  4         �t�bhhK ��h��R�(KK��h�C   5   �   �         �t�bhhK ��h��R�(KK��h�Ch~     �
     M  	      	      	   K   	   �   	   �   	     	   I  	   �  	   U  	   �      �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C!         	         �t�bhhK ��h��R�(KK��h�C T      �  R     +         �t�bhhK ��h��R�(KK��h�C�      �     /      �t�bhhK ��h��R�(KK��h�C1        7  �  r      �t�bhhK ��h��R�(KK
��h�C(   v     
     �   $   o        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C1   #       p     �     �t�bhhK ��h��R�(KK��h�C4   '   -      V   8     �     �   &        �t�bhhK ��h��R�(KK
��h�C(   	      	      	   K   	   U     �t�bhhK ��h��R�(KK��h�C�  q        �t�bhhK ��h��R�(KK��h�C`   �     �
        8     �
     9  V      {  $   �     $   :     �  �        �t�bhhK ��h��R�(KK��h�C;        �t�bhhK ��h��R�(KK��h�C0
      ]  T  '   !      .     �         �t�bhhK ��h��R�(KK	��h�C$      �     �  r  	         �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�CDb  �
     b      s  �
     �   2      2  �               �t�bhhK ��h��R�(KK��h�C M      +   3     4         �t�bhhK ��h��R�(KK��h�C,   {  �          �     �        �t�bhhK ��h��R�(KK��h�C8      -   �  +              <  =           �t�bhhK ��h��R�(KK
��h�C(W   �   t     �  �              �t�bhhK ��h��R�(KK��h�Cd�      
   4  	      	      	   K   	   �   	   I  	   �  	   U  	   /  	   s  	   �     �t�bhhK ��h��R�(KK��h�C    �        8   �        �t�bhhK ��h��R�(KK��h�C4/      -   6        �        >           �t�bhhK ��h��R�(KK��h�C4�  �   +   x      5        `             �t�bhhK ��h��R�(KK��h�C`*      �         D  l        �   f        �      �   ;      0   �     �        �t�bhhK ��h��R�(KK��h�C      2         �        �t�bhhK ��h��R�(KK��h�C u     �  �  �   E        �t�bhhK ��h��R�(KK��h�C,   2   �  Y  ?     2   0   �        �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�C8�      =      [      v    ^   �               �t�bhhK ��h��R�(KK��h�C06  �        F     G     C  /         �t�bhhK ��h��R�(KK��h�CT%   �   .  w  @     
   �        2      �   t     �   �      O        �t�bhhK ��h��R�(KK��h�CH      D  =         �  4      m  >      a      �  �         �t�bhhK ��h��R�(KK��h�C      �            �t�bhhK ��h��R�(KK	��h�C$      A  ?                �t�bhhK ��h��R�(KK��h�CH      c     `   m      /     B  i     %   ^  "   �        �t�bhhK ��h��R�(KK��h�CH      J         )     �   �   S        �     5           �t�bhhK ��h��R�(KK��h�C4     �      5   �      �         C        �t�bhhK ��h��R�(KK��h�C�   -     �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�CT
        2   �   0  p  
   z  �   7      �  �  p  
   z  s   7         �t�bhhK ��h��R�(KK��h�CL@   �   �        /      �  M     {     e     �  g           �t�bhhK ��h��R�(KK��h�CZ   D     �t�bhhK ��h��R�(KK��h�C,�  1        4   �   �      �         �t�bhhK ��h��R�(KK��h�C0]   �     E     F                    �t�bhhK ��h��R�(KK��h�CD   (   H              R  H     4   
   �   �   _         �t�bhhK ��h��R�(KK��h�C4      6  +      �  �        d  G        �t�bhhK ��h��R�(KK��h�Cx     �t�bhhK ��h��R�(KK��h�C�  H     �     �t�bhhK ��h��R�(KK��h�C q               I        �t�bhhK ��h��R�(KK��h�C�   !      �  	         �t�bhhK ��h��R�(KK��h�C0      �     0      k                   �t�bhhK ��h��R�(KK	��h�C$�   �  �  �  �               �t�bhhK ��h��R�(KK��h�C,     1        '   
   �  F         �t�bhhK ��h��R�(KK��h�CD
     (      [      "   >  x      �         0   <         �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C�   J     �t�bhhK ��h��R�(KK��h�C1   #       �        �t�bhhK ��h��R�(KK��h�C8�     K  �     C   �      �     �  �        �t�bhhK ��h��R�(KK��h�Cp�  L  �  M                                      N     O     P  (   N   A     I        �t�bhhK ��h��R�(KK
��h�C(Q  y           �      I         �t�bhhK ��h��R�(KK��h�C<   �      $  �      �  i                       �t�bhhK ��h��R�(KK��h�C8      )   P   ^     �      ^   q   R  F         �t�bhhK ��h��R�(KK��h�C`   �      e     �  i   #  �     !  �  	  S     z     �        �   w         �t�bhhK ��h��R�(KK��h�CP      �     �  5         �           >   a                    �t�bhhK ��h��R�(KK��h�C4
   �     �     F   '      H     �        �t�bhhK ��h��R�(KK��h�C  �   �  �  �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C�   v            �t�bhhK ��h��R�(KK��h�C<M      \  L     
   *         =         �        �t�bhhK ��h��R�(KK��h�C4h  �  O   >   )  C   �  G   |      �         �t�bhhK ��h��R�(KK��h�CT   �            �t�bhhK ��h��R�(KK��h�C47     ;      w   5     �   J   �   8        �t�bhhK ��h��R�(KK	��h�C$T      9        �   �         �t�bhhK ��h��R�(KK��h�C\   �   �  r      �t�bhhK ��h��R�(KK��h�C0         \     (         �           �t�bhhK ��h��R�(KK��h�C@1   #      f        
   3   6     �   �               �t�bhhK ��h��R�(KK��h�C �  T     
     U        �t�bhhK ��h��R�(KK��h�C@   t     /   9   -  (   2   <           �           �t�bhhK ��h��R�(KK	��h�C$                 �         �t�bhhK ��h��R�(KK��h�C<
   V  F         �  �    �     /      {        �t�bhhK ��h��R�(KK��h�C:  �  �   �          �t�bhhK ��h��R�(KK��h�C�        �t�bhhK ��h��R�(KK��h�C�             �t�bhhK ��h��R�(KK��h�C`"   W       X    p      Y  �  h   �     �          Z     [     \        �t�bhhK ��h��R�(KK��h�C\]     �  ^        �         �         _        :      S   Y      Q         �t�bhhK ��h��R�(KK��h�CD*      �  +                   ;  +      `  <        �t�bhhK ��h��R�(KK��h�CD   '   �  �     �  
   a                            �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C<      �   %   �                 k               �t�bhhK ��h��R�(KK��h�CP
   3   6   7  }     o   ?      !      \   2   |     o               �t�bhhK ��h��R�(KK��h�C0   b  �  5         �        Z        �t�bhhK ��h��R�(KK��h�Cc     �t�bhhK ��h��R�(KK��h�C  
         �t�bhhK ��h��R�(KK��h�CD-     b        S  u  �     �     l      �  b        �t�bhhK ��h��R�(KK	��h�C$p      :          �        �t�bhhK ��h��R�(KK��h�C0�  ;  d        <                    �t�bhhK ��h��R�(KK��h�C@�   q   7  &   I     �  �  }     C  �             �t�bhhK ��h��R�(KK��h�C<   d  �     �  �     ~     l      5            �t�bhhK ��h��R�(KK��h�C<      M   �   �         �           <           �t�bhhK ��h��R�(KK��h�C1   #          �t�bhhK ��h��R�(KK��h�C�     �   e           �t�bhhK ��h��R�(KK
��h�C(,   �          	      	         �t�bhhK ��h��R�(KK��h�CD$   �     T           �           �   o               �t�bhhK ��h��R�(KK��h�C<      
   _          |  �     7  J          �t�bhhK ��h��R�(KK��h�C         e  
   c        �t�bhhK ��h��R�(KK	��h�C$�       ^     B   �        �t�bhhK ��h��R�(KK
��h�C(   (   �  �          �        �t�bhhK ��h��R�(KK��h�Cf  �   �   �         �t�bhhK ��h��R�(KK
��h�C(     �           ;   g        �t�bhhK ��h��R�(KK��h�C   J  C      !     �t�bhhK ��h��R�(KK��h�Ch  �     $   �         �t�bhhK ��h��R�(KK	��h�C$#   !   ?      
   �   F         �t�bhhK ��h��R�(KK��h�C=  	         �t�bhhK ��h��R�(KK��h�C�        o  <     �t�bhhK ��h��R�(KK��h�C<"   e   �
     �           /      ^  z           �t�bhhK ��h��R�(KK	��h�C$      3  �     k            �t�bhhK ��h��R�(KK��h�C   4  '   �   i        �t�bhhK ��h��R�(KK��h�C,%   �     j  :   @      X   �        �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6   k        �t�bhhK ��h��R�(KK��h�C8      �  c   �            l     
            �t�bhhK ��h��R�(KK��h�CL   ?   m  *      �  "  n  o  "     u  �         p           �t�bhhK ��h��R�(KK	��h�C$H  �  +            q        �t�bhhK ��h��R�(KK��h�C8%   >  r     �   �            s               �t�bhhK ��h��R�(KK��h�C<            z   
   ,            �  
            �t�bhhK ��h��R�(KK��h�C0v  �        .   s     t              �t�bhhK ��h��R�(KK��h�C0w     ;     u          "   5        �t�bhhK ��h��R�(KK��h�CD*            k         �   Q  R      �     .   �        �t�bhhK ��h��R�(KK��h�CK         Z   �     �t�bhhK ��h��R�(KK��h�C   k  j     /        �t�bhhK ��h��R�(KK��h�CX         8        �   O      ~               0   4   
   _      �        �t�bhhK ��h��R�(KK
��h�C(      )   M   +                 �t�bhhK ��h��R�(KK��h�C@a           �  	      	      	   K   	   U  	   /     �t�bhhK ��h��R�(KK��h�CP   n      �t�bhhK ��h��R�(KK��h�Cv  M             �t�bhhK ��h��R�(KK��h�C0�   7  (   �       .      �   ?         �t�bhhK ��h��R�(KK��h�C   =      �      �t�bhhK ��h��R�(KK��h�C4   (   #   !      �     $   x  
           �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0  �      �  �   �        O  �        �t�bhhK ��h��R�(KK$��h�C�*   H     w     �  �   
   $   E         
   _      �          K       x     `         �     �   �      �  �        �t�bhhK ��h��R�(KK��h�C8V                 �     $  �              �t�bhhK ��h��R�(KK��h�Cq     �t�bhhK ��h��R�(KK��h�CT   �  �  �  �  �  h      �   L     �          v  ;      y        �t�bhhK ��h��R�(KK��h�C       z   ,               �t�bhhK ��h��R�(KK��h�C8T   �                                    �t�bhhK ��h��R�(KK��h�C   �     8   �        �t�bhhK ��h��R�(KK��h�C4
     �      u   p        �   
           �t�bhhK ��h��R�(KK��h�Cg  �           e      �t�bhhK ��h��R�(KK��h�CG     u        �t�bhhK ��h��R�(KK
��h�C(   �  &   `     �  �  �        �t�bhhK ��h��R�(KK��h�C,Z      �               �            �t�bhhK ��h��R�(KK��h�CH^  u            Y  �  :   �   �   Q      �   O  
   �        �t�bhhK ��h��R�(KK��h�C,      �  �  0  �        z        �t�bhhK ��h��R�(KK��h�Ch{        Y           �            �       �      �      �  �      h     �         �t�bhhK ��h��R�(KK��h�CT|           �     I   /   �           ;      }        �           �t�bhhK ��h��R�(KK��h�C     	      	         �t�bhhK ��h��R�(KK��h�C<�      �  �     R            �     v   �        �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK
��h�C(~    @  '   9     ]          �t�bhhK ��h��R�(KK��h�C@"   �           e      @         z   h   H   �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C      �   f     �t�bhhK ��h��R�(KK��h�C,:  
      �     M     {  7         �t�bhhK ��h��R�(KK��h�CP   �      $     �  �   Y  +      �  +      �      U      �        �t�bhhK ��h��R�(KK��h�C!  �     0   <         �t�bhhK ��h��R�(KK��h�C8            �     "     ]  �     Z        �t�bhhK ��h��R�(KK��h�Cp         �   �  �  
   #           �          $  %     >      v            �            �t�bhhK ��h��R�(KK��h�CP      &        �  �   �     '  �     �  �  
         �        �t�bhhK ��h��R�(KK��h�C<   i  �  R         /   9     7         �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C,.  M        
        �            �t�bhhK ��h��R�(KK��h�CD            �     M   T   �   �           i           �t�bhhK ��h��R�(KK��h�C         �           �t�bhhK ��h��R�(KK��h�C   �      �t�bhhK ��h��R�(KK��h�C<�  N  
   8     ^   &  �     
      �  �        �t�bhhK ��h��R�(KK��h�C   �  
   �     �t�bhhK ��h��R�(KK��h�C<      5  �      \   �        &     
   U        �t�bhhK ��h��R�(KK��h�C              �t�bhhK ��h��R�(KK��h�Cq            �t�bhhK ��h��R�(KK��h�C\
   3   6   �  ?      !      #        �      $   �  �  �      �     �         �t�bhhK ��h��R�(KK��h�C0   >   �       �   *   �  �  V         �t�bhhK ��h��R�(KK��h�C4�  9     W     (           )  �
        �t�bhhK ��h��R�(KK��h�C@�     �           �
  :   �  
   _      �  �        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�CD      P           *         E  �        �   �         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C1   #       +        �t�bhhK ��h��R�(KK��h�Ct   $   V  �     �     C   w         A              
      A     Z        �         �        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C �        	      	         �t�bhhK ��h��R�(KK��h�C8   �     �      *  L     �         �        �t�bhhK ��h��R�(KK��h�C4#   !      �        (      ^   Q           �t�bhhK ��h��R�(KK/��h�C�   R  %     �                             �  u      �     �     A   �     X         J   a   !         .   �      �     {      _     B     �  �         �t�bhhK ��h��R�(KK��h�Cd         0   �     �  �        (   �     �      �     w   �   �      `   /         �t�bhhK ��h��R�(KK��h�C4   W     :   �  �  �        ^            �t�bhhK ��h��R�(KK��h�C4�   ,   9  �     �      �  )      u         �t�bhhK ��h��R�(KK��h�CP        �   f     �         1   #   
   3   6     �   �            �t�bhhK ��h��R�(KK��h�C!      ,         �t�bhhK ��h��R�(KK��h�C0
        �     e  �                 �t�bhhK ��h��R�(KK��h�C�              �t�bhhK ��h��R�(KK��h�Cl�     �     +  �        �                       �      �     +  �     �   �         �t�bhhK ��h��R�(KK��h�C@,  L  �            �  &      H  �    
   �        �t�bhhK ��h��R�(KK��h�C>   �   v   r      �t�bhhK ��h��R�(KK��h�C,      )   b      #   !      �        �t�bhhK ��h��R�(KK��h�C          	      	         �t�bhhK ��h��R�(KK��h�Cb      x   
   �     �t�bhhK ��h��R�(KK	��h�C$`   b           �  �        �t�bhhK ��h��R�(KK��h�CW      �t�bhhK ��h��R�(KK��h�C    W  �   '      e         �t�bhhK ��h��R�(KK��h�CL2      =      �     �     �  �   �  7      �     J  /         �t�bhhK ��h��R�(KK��h�C0�        -  p         �      �        �t�bhhK ��h��R�(KK��h�C�     A   �     �t�bhhK ��h��R�(KK��h�C4Z         �     �  �      �     �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C8
   �   F   ?      -   1     \        +        �t�bhhK ��h��R�(KK��h�C0o  �      /      �      	      	         �t�bhhK ��h��R�(KK��h�C5     �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK	��h�C$�        .                 �t�bhhK ��h��R�(KK��h�C4*      �   F  &      U        8   �        �t�bhhK ��h��R�(KK��h�C      	      	   K      �t�bhhK ��h��R�(KK��h�Cp   �   :      Q   �  Y   �   Q     a   ;      f      �   �        .   %   �          f        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C 1   #       �              �t�bhhK ��h��R�(KK��h�C[      �     �t�bhhK ��h��R�(KK��h�C8                         <               �t�bhhK ��h��R�(KK
��h�C(�      �  	      	   K   	   �      �t�bhhK ��h��R�(KK��h�C%   �  O     �t�bhhK ��h��R�(KK
��h�C(         '  �  �   B   �        �t�bhhK ��h��R�(KK��h�C�      	      	         �t�bhhK ��h��R�(KK��h�C0�  �  .        5      �  
   6        �t�bhhK ��h��R�(KK��h�C/  q   0         �t�bhhK ��h��R�(KK��h�Cd�  �   |      �      �     �        1     �            J   �     �     W         �t�bhhK ��h��R�(KK��h�Cd      J   a   �  �       y              c  p            =      �     �         �t�bhhK ��h��R�(KK��h�Cd-      �     �     2   (   /         �  �  �   �      2   5   [         !  #        �t�bhhK ��h��R�(KK��h�C`      0   [                        ~            :     �     "              �t�bhhK ��h��R�(KK��h�C,b   #   "      �  V      J   z         �t�bhhK ��h��R�(KK��h�C2  R      �        �t�bhhK ��h��R�(KK��h�CT         �  G      �        =      [      C     "   $   �   �        �t�bhhK ��h��R�(KK��h�Cp9   �  (         j  <         �  �   |     x      "   >  D     �   �  V   2      0   <         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C0   Y      O   5      7                 �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK	��h�C$#     �   z      c  X  r      �t�bhhK ��h��R�(KK��h�C�   �     �     �t�bhhK ��h��R�(KK��h�C4V     3  &   N   
   ,                     �t�bhhK ��h��R�(KK��h�C1   #       	  l         �t�bhhK ��h��R�(KK��h�C          I   �  C         �t�bhhK ��h��R�(KK
��h�C(   E  j        k  j  /        �t�bhhK ��h��R�(KK��h�C<      b   "   W  W      �  \         0           �t�bhhK ��h��R�(KK��h�C,�     S     '   
   �   B   }         �t�bhhK ��h��R�(KK��h�C8   �  �     �   �  �  �  �  �  0  ;        �t�bhhK ��h��R�(KK
��h�C(�     I     �        �         �t�bhhK ��h��R�(KK��h�CL�      \  �   �      4     
   F  F      �   �  $     �        �t�bhhK ��h��R�(KK��h�C�     �  	         �t�bhhK ��h��R�(KK��h�Cl�   &   �     �      G       %   H  �     �   "   �  �  �  �   �     Y  �      �        �t�bhhK ��h��R�(KK��h�CD      �                    �  �          �        �t�bhhK ��h��R�(KK��h�C8?         �  �   I  V         =      n         �t�bhhK ��h��R�(KK��h�C�     A   �      �t�bhhK ��h��R�(KK��h�C 1   #   
   3   6   t        �t�bhhK ��h��R�(KK��h�C�  4   �     �t�bhhK ��h��R�(KK��h�C1   #       i        �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C�  5     �t�bhhK ��h��R�(KK��h�C4   &   a      +   J  
   �   $     k        �t�bhhK ��h��R�(KK	��h�C$6  �           �           �t�bhhK ��h��R�(KK��h�C�           �t�bhhK ��h��R�(KK��h�C7  �  
   �     �t�bhhK ��h��R�(KK��h�C0      �   �         )  +   
   &        �t�bhhK ��h��R�(KK��h�C4      6  +      �  �        d  G        �t�bhhK ��h��R�(KK��h�Cd      V  �  �        5   [         U   @     �     e      �      �      �        �t�bhhK ��h��R�(KK��h�C`      D   &   D  0   4   >   P  �   �  �        N   �        .   �     �        �t�bhhK ��h��R�(KK��h�CH      �     o  ~             ?      8  
   8           �t�bhhK ��h��R�(KK��h�CZ      �            �t�bhhK ��h��R�(KK��h�C�  R      �t�bhhK ��h��R�(KK��h�C,   �                            �t�bhhK ��h��R�(KK��h�C4�  �          �        �        �     �t�bhhK ��h��R�(KK��h�C   �  
   �     �t�bhhK ��h��R�(KK��h�C[   "   �     �t�bhhK ��h��R�(KK��h�C�      D      �t�bhhK ��h��R�(KK��h�C�     �     �t�bhhK ��h��R�(KK��h�C@      ]  �     �  Q     �  &   �   �             �t�bhhK ��h��R�(KK��h�C0   �  I   �     Y      O   �  �         �t�bhhK ��h��R�(KK
��h�C(1   #   
   3   6   �     �        �t�bhhK ��h��R�(KK��h�C@   &   T   �     E       	     �           
        �t�bhhK ��h��R�(KK��h�C@�     �      N   �     �   �     %   �      I         �t�bhhK ��h��R�(KK��h�C0�   �     �   9  �     �  i   �         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK	��h�C$~     l      :        �     �t�bhhK ��h��R�(KK��h�C E      �  	      	         �t�bhhK ��h��R�(KK��h�C   
   �     �t�bhhK ��h��R�(KK��h�C
      5     �        �t�bhhK ��h��R�(KK��h�C<
   �   F   ?      �     �     #   !      P        �t�bhhK ��h��R�(KK��h�C4   .   (   �     a   �   <       <        �t�bhhK ��h��R�(KK��h�C8�
     )   N      �
                 �        �t�bhhK ��h��R�(KK��h�C<�   �        >   ;  �       %   &             �t�bhhK ��h��R�(KK��h�C0d  
   \   8   �  �  �  �     �        �t�bhhK ��h��R�(KK��h�CL
   Z        R  �     �          �     	     �   S         �t�bhhK ��h��R�(KK��h�CJ     /      �t�bhhK ��h��R�(KK��h�C    �  �   0  B   [        �t�bhhK ��h��R�(KK
��h�C(�  a  �     �  9   �  �        �t�bhhK ��h��R�(KK��h�C@      �  #      S     �  
   3   6   �             �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C`   �           %                    �
     8   �     $   A     $   p         �t�bhhK ��h��R�(KK��h�CT�        �  �            �  K  G   /      T  �   D   %   �  	        �t�bhhK ��h��R�(KK��h�C0  �     >     U     �   �   B         �t�bhhK ��h��R�(KK��h�C4   (   #   !      �     $   x  
   k        �t�bhhK ��h��R�(KK��h�C@a     G  P     $   �   �  s   �   y      �   <        �t�bhhK ��h��R�(KK��h�C�  �      �t�bhhK ��h��R�(KK��h�C@k     e      �  �     �     �   
   H   B           �t�bhhK ��h��R�(KK��h�C	  �     �  �  �     �t�bhhK ��h��R�(KK��h�C   (   �  9   �        �t�bhhK ��h��R�(KK��h�C      @          �t�bhhK ��h��R�(KK��h�C�  �          �     �t�bhhK ��h��R�(KK��h�C01   #   
   3   6   �     �     �        �t�bhhK ��h��R�(KK(��h�C��           P     2      �            �      �     �     =  i   A      .   
   _      L  �     >     �          X     d        �t�bhhK ��h��R�(KK��h�C8�  	  �   	  9   �            �
              �t�bhhK ��h��R�(KK��h�Cx   D         �     �   S        #     D      �   �           V     �      �   	  V              �t�bhhK ��h��R�(KK��h�C\               k         &        W   �  $   ;         �        �        �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C4      �  
         �  )   
   A   }         �t�bhhK ��h��R�(KK��h�Ce         �t�bhhK ��h��R�(KK
��h�C(#   !   '   
   �   �  ?  F         �t�bhhK ��h��R�(KK��h�C<�      �  v   �        �     ,      $   @        �t�bhhK ��h��R�(KK��h�C�      /              �t�bhhK ��h��R�(KK��h�C0      �      A     �   �     "        �t�bhhK ��h��R�(KK��h�C8�  	  +            �     �         �        �t�bhhK ��h��R�(KK��h�CL      q   B  �     �     ,        �  �  C  �     �        �t�bhhK ��h��R�(KK��h�CD   (   z         A     _  *      a          �
        �t�bhhK ��h��R�(KK��h�CX      -   P   n   ^   %  �  	     �     �  	     �                    �t�bhhK ��h��R�(KK��h�C0�        �  �            ;   �        �t�bhhK ��h��R�(KK��h�C4   5   &        �      		     $   �         �t�bhhK ��h��R�(KK��h�C,D        �           �            �t�bhhK ��h��R�(KK��h�CH*         E  H        ;      G        �  $   E   �        �t�bhhK ��h��R�(KK��h�C4�     T   a   e  �     l  �     D         �t�bhhK ��h��R�(KK��h�CH   `   b  �   �     e  9   y     &      
     �          �t�bhhK ��h��R�(KK��h�CB  �     �  �        �t�bhhK ��h��R�(KK��h�C@         �      �      7      �  F     +  �        �t�bhhK ��h��R�(KK��h�C   �  �             �t�bhhK ��h��R�(KK��h�Cd\      j     	      	      	   K   	   �   	   �   	     	   �   	   �  	   �  	   /     �t�bhhK ��h��R�(KK��h�C4E   &   �  y         �  �   �   s   7         �t�bhhK ��h��R�(KK��h�C,�     \   �         �     :        �t�bhhK ��h��R�(KK��h�C�   ]  �               �t�bhhK ��h��R�(KK��h�C   �              �t�bhhK ��h��R�(KK��h�C
	  =     �     �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C,^   �   �  �     R      �   �         �t�bhhK ��h��R�(KK��h�C@�      (  �  u      �      ,   �                    �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C4]   P        �                 G        �t�bhhK ��h��R�(KK��h�C8#   !      �  '   
   3   6   �  t              �t�bhhK ��h��R�(KK��h�C\      r  '  (      !      p      ,                  p      R      X         �t�bhhK ��h��R�(KK��h�C �     m  �                �t�bhhK ��h��R�(KK��h�C,m  �  �     �           X        �t�bhhK ��h��R�(KK��h�C<1   #      ,   �       �  
   3   6   	  �         �t�bhhK ��h��R�(KK��h�Cd   �      $     �  �   Y  +      �  +      �            U      �     	           �t�bhhK ��h��R�(KK
��h�C(   '      �     	     H        �t�bhhK ��h��R�(KK��h�C0�        �     y     �      �        �t�bhhK ��h��R�(KK��h�C�   p      �t�bhhK ��h��R�(KK��h�CI               �t�bhhK ��h��R�(KK��h�C0      h  �  �  �     S      5        �t�bhhK ��h��R�(KK��h�C,*        �  &      �     E          �t�bhhK ��h��R�(KK��h�CP�          �                 W       b  �      �  	        �t�bhhK ��h��R�(KK��h�C	  J  
            �t�bhhK ��h��R�(KK��h�C K     	                 �t�bhhK ��h��R�(KK��h�C	     �      �         �t�bhhK ��h��R�(KK
��h�C(         L  +         �        �t�bhhK ��h��R�(KK��h�C,-   n  �  7      :   M     @         �t�bhhK ��h��R�(KK��h�CH�   =  �  >     ,      A   �         E  9      �            �t�bhhK ��h��R�(KK��h�CP   @   '      -   �   e     �   
   �        /     �      K         �t�bhhK ��h��R�(KK��h�CX:   Q     z  (      M      +      j  �     �   �
     �     �  �
        �t�bhhK ��h��R�(KK��h�CP)   A   6        �            4   
   _      X  �     R  4         �t�bhhK ��h��R�(KK��h�C�  �     %   �         �t�bhhK ��h��R�(KK��h�C   +     �t�bhhK ��h��R�(KK��h�C�  
   ,      �t�bhhK ��h��R�(KK��h�C8     
   \   �             Y              �t�bhhK ��h��R�(KK
��h�C(�  �           M     	        �t�bhhK ��h��R�(KK��h�C,f         �  h        g            �t�bhhK ��h��R�(KK��h�CP      R  H           �          �   �     8   E  
   _         �t�bhhK ��h��R�(KK��h�C,j   �    �   �     �  
   �  N     �t�bhhK ��h��R�(KK��h�C,E      f   O  (  �      �  E         �t�bhhK ��h��R�(KK��h�CL�   v              �  $   k            �   s   7               �t�bhhK ��h��R�(KK	��h�C$�  (   �                    �t�bhhK ��h��R�(KK��h�C4         �  +      �     �  $           �t�bhhK ��h��R�(KK��h�C	  	         �t�bhhK ��h��R�(KK��h�C)     �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�Cl         .         D   ~   G      �  �           A   �  �
  �     �   f   Z  9            �t�bhhK ��h��R�(KK��h�CPB   P          �     �     �     �           	     �        �t�bhhK ��h��R�(KK��h�CD              �           (      v     �           �t�bhhK ��h��R�(KK��h�C\y      �  $   �     1   Q  S     d  
            �  �      R  g         �t�bhhK ��h��R�(KK��h�C        �  �        �t�bhhK ��h��R�(KK	��h�C$/   9   �  7   5      �
        �t�bhhK ��h��R�(KK��h�C             �t�bhhK ��h��R�(KK��h�C�     S  �     �t�bhhK ��h��R�(KK��h�CH   <               *  3   �  
   A   _     �  B            �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C0!      .  '   
   T     u      X         �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C@   �     �t�bhhK ��h��R�(KK��h�C�  �      N      .      �t�bhhK ��h��R�(KK��h�CD   �   �     	  	        v  �  �  u  c   �           �t�bhhK ��h��R�(KK��h�CP.  "   �     �          <     �     /     ~   �               �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�C8   @   '   H   �   	     )   �   �      /         �t�bhhK ��h��R�(KK��h�C8               �  6     �     8   �        �t�bhhK ��h��R�(KK��h�CP1   #      �             �   f  
   3   6     �   �               �t�bhhK ��h��R�(KK��h�C   y     �t�bhhK ��h��R�(KK��h�C�   	  	         �t�bhhK ��h��R�(KK��h�C�  Y  �         �t�bhhK ��h��R�(KK��h�Cl     �  Q  p      u      �     �     �   �  �     A        �        z   "           �t�bhhK ��h��R�(KK��h�C<
   3   6   �     j   4   '      #   !      �        �t�bhhK ��h��R�(KK��h�CL      0   [         
   _      8   �     $   \  5   0  <         �t�bhhK ��h��R�(KK��h�CR      T     �t�bhhK ��h��R�(KK��h�C�   =     �t�bhhK ��h��R�(KK��h�CL              /               b   x   "                     �t�bhhK ��h��R�(KK��h�C�  �     �t�bhhK ��h��R�(KK��h�C       �  �   7  �        �t�bhhK ��h��R�(KK��h�Cm      �         :     �t�bhhK ��h��R�(KK��h�C
   �  �  [  �        �t�bhhK ��h��R�(KK��h�C<N  7  P   �  :      	      	      	   K   	   �      �t�bhhK ��h��R�(KK��h�C	  �     �t�bhhK ��h��R�(KK��h�C@7         !  �     @      4        n  U  o        �t�bhhK ��h��R�(KK��h�Ch      \  	           �  c         ]     (        ^  )      $   k         X         �t�bhhK ��h��R�(KK��h�CH   &   �  "   �        	  u     �   "   q   �     u        �t�bhhK ��h��R�(KK��h�C`      �                  V     �          �                     �         �t�bhhK ��h��R�(KK��h�CK         �      �     �t�bhhK ��h��R�(KK��h�C�     x  �           �t�bhhK ��h��R�(KK	��h�C$�      �   9   z  q   .        �t�bhhK ��h��R�(KK��h�C O     	  �      ?        �t�bhhK ��h��R�(KK
��h�C(            �        N  �     �t�bhhK ��h��R�(KK��h�C,_        �  �     �      �        �t�bhhK ��h��R�(KK��h�C4     G  �   [      �      G     �        �t�bhhK ��h��R�(KK��h�C[      �      �t�bhhK ��h��R�(KK��h�C8   (   !      \      ]  �  
   3   6   	        �t�bhhK ��h��R�(KK��h�C�   >   5  �        �t�bhhK ��h��R�(KK��h�C !      �  	      	         �t�bhhK ��h��R�(KK��h�CHk  �  	  
   N              V  �      O     9           �t�bhhK ��h��R�(KK��h�C   �  	      	         �t�bhhK ��h��R�(KK��h�C	  �          �t�bhhK ��h��R�(KK��h�C8
   �     5     -   \   '     $   E   W        �t�bhhK ��h��R�(KK��h�C<         .   �     �  >      w   v   �           �t�bhhK ��h��R�(KK��h�C8      '   P  �     �        �              �t�bhhK ��h��R�(KK��h�C,     &      �         �   	  r      �t�bhhK ��h��R�(KK��h�C X     �  
   ]  L         �t�bhhK ��h��R�(KK��h�C1   #       �  4         �t�bhhK ��h��R�(KK��h�C@   �                  �     Q     �  �  �        �t�bhhK ��h��R�(KK��h�C0b     �     =  �  >         �        �t�bhhK ��h��R�(KK��h�C    E  j     j  /        �t�bhhK ��h��R�(KK��h�C4*   r  $  �     0     D     +  2        �t�bhhK ��h��R�(KK	��h�C$   �  +  '   �  �           �t�bhhK ��h��R�(KK��h�C#  �     p  r      �t�bhhK ��h��R�(KK
��h�C(�     !	     -      P           �t�bhhK ��h��R�(KK��h�C"	  �     �t�bhhK ��h��R�(KK��h�Cl�   q   7  &   �  Y  �   �           �   O      +  l           q     +   '      �        �t�bhhK ��h��R�(KK��h�C02      �   �   >  �  y                  �t�bhhK ��h��R�(KK��h�C<      '   H   �     �             #	           �t�bhhK ��h��R�(KK��h�C�  	         �t�bhhK ��h��R�(KK	��h�C$   @   '   �       `        �t�bhhK ��h��R�(KK��h�C@$	  �         �      �  �        �  �     `        �t�bhhK ��h��R�(KK��h�C8�   ^                        �     Y        �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6   �  t              �t�bhhK ��h��R�(KK��h�C4*   �     a     2   =      Z     �        �t�bhhK ��h��R�(KK	��h�C$     �  Y  �      7         �t�bhhK ��h��R�(KK��h�C<
   �   F   ?      �     �     #   !      P        �t�bhhK ��h��R�(KK��h�C\   f   s  �      2   [  :   %	        '   �  �          d   b  (  ]         �t�bhhK ��h��R�(KK��h�C <         0   �  
   �      �t�bhhK ��h��R�(KK��h�CD1   #      b     ,     �   p   
   3   6   �     /         �t�bhhK ��h��R�(KK��h�C2   >   2     �        �t�bhhK ��h��R�(KK
��h�C(   >   =      \  �  :   W         �t�bhhK ��h��R�(KK
��h�C(q     �     �  	      	         �t�bhhK ��h��R�(KK��h�CH�     )   �     �  �     \   �  &         �
    ]        �t�bhhK ��h��R�(KK*��h�C�         O         Y      Q      �     x     J   �                �        .   
   �     
               \  �     5      7  L        �t�bhhK ��h��R�(KK��h�C1   #               �t�bhhK ��h��R�(KK��h�C0            �     �        K        �t�bhhK ��h��R�(KK��h�C        �t�bhhK ��h��R�(KK��h�C�
  	      	         �t�bhhK ��h��R�(KK��h�CL      ,  %   �                    k      l                 �t�bhhK ��h��R�(KK��h�Cd      -   �  �      �   �     �  �  '  G   C         &	     �     8   �   S        �t�bhhK ��h��R�(KK��h�C8      -   �  ^  
        "   �     �        �t�bhhK ��h��R�(KK��h�C �      '	        	         �t�bhhK ��h��R�(KK
��h�C(�     �        �  �  �        �t�bhhK ��h��R�(KK
��h�C(!         N  �  	      	         �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�CtY      �       X     -  J  C      �   h   �  �     X     �     �  �      (	     Y      �     �t�bhhK ��h��R�(KK��h�C8)   �  �  =     %      �   �  i   A   =        �t�bhhK ��h��R�(KK��h�C4        J  �     K     X               �t�bhhK ��h��R�(KK��h�C    (   [      �            �t�bhhK ��h��R�(KK��h�C4[      C     	      	      	   �  	   �      �t�bhhK ��h��R�(KK��h�C,N     �      d      	      	         �t�bhhK ��h��R�(KK��h�C   �  g   �            �t�bhhK ��h��R�(KK��h�C@              0   L   G      �  Z        J         �t�bhhK ��h��R�(KK
��h�C($  �  �   .        O  �        �t�bhhK ��h��R�(KK��h�C      �  �        �t�bhhK ��h��R�(KK��h�C`   `   �            .   Y  �  i   s   7      &   �  �  �  �      �      �        �t�bhhK ��h��R�(KK
��h�C(�    
         $   �            �t�bhhK ��h��R�(KK��h�C,      B   �     �  	      	         �t�bhhK ��h��R�(KK��h�C|      �      R          /  �       �     �      -  �     _     �        �     /   �   )	        �t�bhhK ��h��R�(KK��h�C4             0                       �t�bhhK ��h��R�(KK��h�CLq   �  �  �         �  x                 *   �   
  4         �t�bhhK ��h��R�(KK��h�CP      �        /  i        f   ?     /  i  �  +               �t�bhhK ��h��R�(KK��h�Cb   #   G   W         �t�bhhK ��h��R�(KK��h�CH*      �         �     C  W            ;      �   �        �t�bhhK ��h��R�(KK
��h�C(      c     +     �  �         �t�bhhK ��h��R�(KK��h�C?      �     �        �t�bhhK ��h��R�(KK
��h�C(      -   P         �  *	        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C4   (   1     \   ]   /  8   @     �        �t�bhhK ��h��R�(KK��h�C4   �        `  N               a        �t�bhhK ��h��R�(KK��h�C8#   !         =      �   ?      
   �  F         �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C,      �   >      a      �          �t�bhhK ��h��R�(KK��h�C8   &   =      �  4   y   8   3  4     c         �t�bhhK ��h��R�(KK��h�C �   �  ^   �  �           �t�bhhK ��h��R�(KK��h�C<1   #         U        
   3   6   �
              �t�bhhK ��h��R�(KK��h�C<   X   '   )               �   p      B            �t�bhhK ��h��R�(KK��h�C4�     �  �      ,      A   �      �        �t�bhhK ��h��R�(KK��h�C E         	      	         �t�bhhK ��h��R�(KK��h�CH   .   W      b     �     �     f   �      &     �        �t�bhhK ��h��R�(KK��h�C,Y      O   &   -   F  C   
   H        �t�bhhK ��h��R�(KK��h�CS            �t�b�
0      hhK ��h��R�(KK��h�CT         m      �     A   �     +	        M   �      �              �t�bhhK ��h��R�(KK��h�CP        i          $   n            �             ]         �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK��h�C   x         �t�bhhK ��h��R�(KK��h�C    	      	      	   K      �t�bhhK ��h��R�(KK��h�C�  	      	         �t�bhhK ��h��R�(KK��h�Cd      "        s  �   [  :   %	           '   �  �          d   b  (  ]         �t�bhhK ��h��R�(KK��h�CD%     m  �            �  c           �     u         �t�bhhK ��h��R�(KK��h�C,      N   :      �     �   �         �t�bhhK ��h��R�(KK��h�CX!               	      	   K   	   �   	   I  	   U  	   /  	   �  	   �     �t�bhhK ��h��R�(KK��h�CdT      d     (   �      �   �   �     d  �   �  
   _      L  �     d     �        �t�bhhK ��h��R�(KK��h�CD$  �  �  �     >   �  $   0     *  �   �     �        �t�bhhK ��h��R�(KK��h�C0I   u      ;      0   �   !               �t�bhhK ��h��R�(KK��h�C  p      u      �t�bhhK ��h��R�(KK��h�CHw  �  (   #   !      ]   �   s     
   �  F         e        �t�bhhK ��h��R�(KK��h�C0�  "        Q     /   9     7         �t�bhhK ��h��R�(KK��h�C,1   #   
   3   6   �     �  �         �t�bhhK ��h��R�(KK��h�C0�  �       6     �     
            �t�bhhK ��h��R�(KK	��h�C$         f     M   ,	        �t�bhhK ��h��R�(KK��h�C0�     2     :     �   +     -	        �t�bhhK ��h��R�(KK��h�CX      '   -   �        �      �        .         M  �        �        �t�bhhK ��h��R�(KK��h�C,�   �   2      T          <        �t�bhhK ��h��R�(KK��h�C C  �     M     {        �t�bhhK ��h��R�(KK��h�C!           �        �t�bhhK ��h��R�(KK��h�CL�  g     �        ;            /      ;      )	  h   �         �t�bhhK ��h��R�(KK��h�Ch      )        <      x   "   Q  	     �           "   <              .            �t�bhhK ��h��R�(KK	��h�C$4   
   A      	      	         �t�bhhK ��h��R�(KK��h�C4      ]  I        �  �   !      �         �t�bhhK ��h��R�(KK��h�C�  �         �t�bhhK ��h��R�(KK��h�C   �               �t�bhhK ��h��R�(KK
��h�C(�     W  .	     N       r      �t�bhhK ��h��R�(KK��h�C      �t�bhhK ��h��R�(KK��h�C4*               :      n         �          �t�bhhK ��h��R�(KK��h�C4!         ?      
   �  F      
            �t�bhhK ��h��R�(KK��h�C@*   h     �  /  `        $   /	     �  b           �t�bhhK ��h��R�(KK��h�CTN  �     �  	      	      	   K   	   �   	     	   �  	   �   	   �     �t�bhhK ��h��R�(KK��h�C@1   #         �  `   �  
   3   6   �  g  �   �        �t�bhhK ��h��R�(KK��h�C<   @   '      �   5     ]     4     �   5        �t�bhhK ��h��R�(KK��h�Cq     �t�bhhK ��h��R�(KK
��h�C(   �           0	  �           �t�bhhK ��h��R�(KK��h�C      1	  2	        �t�bhhK ��h��R�(KK	��h�C$�     I  �     3	           �t�bhhK ��h��R�(KK	��h�C$T      D   4	  �  �   �        �t�bhhK ��h��R�(KK��h�C   �  �         �t�bhhK ��h��R�(KK��h�Ci     �  5	  	         �t�bhhK ��h��R�(KK��h�C�     �  �      �t�bhhK ��h��R�(KK��h�C8   �      �     %   �  6	  7	  �      D         �t�bhhK ��h��R�(KK��h�C,   B        �      �     U        �t�bhhK ��h��R�(KK��h�C   �  T     j        �t�bhhK ��h��R�(KK
��h�C(_        	      	     	   �      �t�bhhK ��h��R�(KK��h�C01   #   
   3   6         �     �         �t�bhhK ��h��R�(KK��h�CZ      �      �     �t�bhhK ��h��R�(KK��h�C   �      �  �     �t�bhhK ��h��R�(KK��h�Ck          1        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C /  ^  @     �  �         �t�bhhK ��h��R�(KK��h�C<   �        
      \        �        ?        �t�bhhK ��h��R�(KK��h�C<�   	  V  �     D   ~   �   e  i   G   �   8        �t�bhhK ��h��R�(KK��h�CK             �     �t�bhhK ��h��R�(KK��h�C4      ,  ?      �  �      �  �  �        �t�bhhK ��h��R�(KK��h�CH      G        j   4         �  �  V     v      	        �t�bhhK ��h��R�(KK	��h�C$#  �   �   �  8	     �        �t�bhhK ��h��R�(KK��h�C8        �  O      �t�bhhK ��h��R�(KK
��h�C(I   k  �  �     �     9	        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C,d  
     �     %        5         �t�bhhK ��h��R�(KK��h�C<#   !         �     (      G         $   k         �t�bhhK ��h��R�(KK��h�C4�  '                L   T   �   �        �t�bhhK ��h��R�(KK��h�C       �   �      I         �t�bhhK ��h��R�(KK��h�C#     �   r      �t�bhhK ��h��R�(KK��h�C{      �t�bhhK ��h��R�(KK��h�CL*         8   �   �      @      &      F  +           <        �t�bhhK ��h��R�(KK��h�CDE   &   r  �      W   �     �  y               �        �t�bhhK ��h��R�(KK��h�Cl  :	     ;	        �t�bhhK ��h��R�(KK��h�C<�     a   
  �     O     %            m        �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C  n  
   4     �t�bhhK ��h��R�(KK��h�C          �      I         �t�bhhK ��h��R�(KK��h�C<            &   r     2  �     �  g   $	        �t�bhhK ��h��R�(KK��h�C  �   m     �        �t�bhhK ��h��R�(KK��h�CX              W  V   X        S   i   ,                 
   �         �t�bhhK ��h��R�(KK��h�CP�      L   G      o           .      m      p     <	              �t�bhhK ��h��R�(KK��h�C@            h  �       �  �     q     �        �t�bhhK ��h��R�(KK��h�C8
      =    +         r  �  	      	         �t�bhhK ��h��R�(KK��h�C\         m      s     �           M   �      �                x          �t�bhhK ��h��R�(KK��h�Ct      �           �        
   _      �        �     �     s        ;         r  �        �t�bhhK ��h��R�(KK��h�C �      d   8  �  �        �t�bhhK ��h��R�(KK��h�C !         	      	         �t�bhhK ��h��R�(KK��h�CP*      �  
   %       &   �                       t  �        �t�bhhK ��h��R�(KK��h�C0   Y     �   '      �     q           �t�bhhK ��h��R�(KK��h�C,  I        	      	   K   	   �      �t�bhhK ��h��R�(KK��h�Cb   #   "   $   �        �t�bhhK ��h��R�(KK��h�C0+     -	  �   +   =	        �  �        �t�bhhK ��h��R�(KK��h�C4     �   �      >	     �         �        �t�bhhK ��h��R�(KK	��h�C$      U     �     ?	        �t�bhhK ��h��R�(KK��h�C !        	      	         �t�bhhK ��h��R�(KK��h�C0   	        �   k     a     �        �t�bhhK ��h��R�(KK��h�C,Z      �               �            �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�C<N  �        ,      	   K   	   �   	     	   �      �t�bhhK ��h��R�(KK��h�C43  �        �     '  
      �   �        �t�bhhK ��h��R�(KK��h�C  (         �        �t�bhhK ��h��R�(KK��h�CD   @	  �
     .      u  �  
               <        �t�bhhK ��h��R�(KK��h�C         b  �           �t�bhhK ��h��R�(KK��h�C,      �      �        �  �         �t�bhhK ��h��R�(KK��h�C4      �        0        �             �t�bhhK ��h��R�(KK��h�C,           T   A	  2   v           �t�bhhK ��h��R�(KK��h�CDM     
               �   A   w        D  v   �        �t�bhhK ��h��R�(KK1��h�CĦ     N   �     .   *   2      :      Q         S         m   
   �     x  �   �        m      �        �  �      x     �     �   F     *   �     
   A           �t�bhhK ��h��R�(KK
��h�C(#   !   ?      
   @   �   F         �t�bhhK ��h��R�(KK��h�C<^   �                  P   !   �   B	     �        �t�bhhK ��h��R�(KK��h�CH   @      �  u   ;      0   �     y  �   h   %   �           �t�bhhK ��h��R�(KK��h�C0W  �     �  B  8   �        t        �t�bhhK ��h��R�(KK��h�C    4  
   t         �t�bhhK ��h��R�(KK��h�C0      0   �     C	     $   �   �        �t�bhhK ��h��R�(KK��h�CZ   .     z        �t�bhhK ��h��R�(KK��h�C   	      	         �t�bhhK ��h��R�(KK��h�CLD   (   �  �  {   �       �              �  �      �        �t�bhhK ��h��R�(KK��h�C         �t�bhhK ��h��R�(KK��h�C         {         �t�bhhK ��h��R�(KK��h�C +     )   �     �        �t�bhhK ��h��R�(KK��h�C�     �t�bhhK ��h��R�(KK��h�C@\      �      �     M    
        Q      ~         �t�bhhK ��h��R�(KK��h�C 5   �      �      �  r      �t�bhhK ��h��R�(KK��h�C0R      ]           S                  �t�bhhK ��h��R�(KK	��h�C$      2     c  X           �t�bhhK ��h��R�(KK��h�CL  h   �  �   :      B   ?     X     ,         �     a   �     �t�bhhK ��h��R�(KK��h�CX   5  _  D   �     �   f     _  C      ,   �              �  �        �t�bhhK ��h��R�(KK��h�Ch   D	  
   �         �  ?               ^   %        �  ?     �   �  �  
   T        �t�bhhK ��h��R�(KK��h�C�      D      V     �t�bhhK ��h��R�(KK��h�CN  7      �t�bhhK ��h��R�(KK��h�CD-   H   �    �   �      .      �     !       @        �t�bhhK ��h��R�(KK��h�CL         8   �   �           &      F  +           <        �t�bhhK ��h��R�(KK
��h�C(�  {           �             �t�bhhK ��h��R�(KK��h�C   �     �t�bhhK ��h��R�(KK��h�CX   >   =         �  4   
   _      {   y   8   4         P   {     c         �t�bhhK ��h��R�(KK��h�CX"   X   E	     g           2      .   �  �     |     F	  �     }        �t�bhhK ��h��R�(KK��h�Cp            Z        S   Y      Q      Q     Q         x        ;      y  ^              �t�bhhK ��h��R�(KK	��h�C$"   G	        )   �   +        �t�bhhK ��h��R�(KK��h�CX     �   �     �t�bhhK ��h��R�(KK��h�C�  T     �t�bhhK ��h��R�(KK��h�Cb      	      	         �t�bhhK ��h��R�(KK��h�C<�   7        ;      �  e  ,                     �t�bhhK ��h��R�(KK��h�C,f   �     @        �  
   ~        �t�bhhK ��h��R�(KK��h�C )     T      $   �        �t�bhhK ��h��R�(KK��h�C     �t�bhhK ��h��R�(KK��h�C,   �   �             G   �         �t�bhhK ��h��R�(KK��h�Cp   Y        S   X  i   ,            �  �  �     T        �  P        �                �t�bhhK ��h��R�(KK��h�CP   R      �t�bhhK ��h��R�(KK��h�C0      :     �   
   ,      
            �t�bhhK ��h��R�(KK��h�C          �t�bhhK ��h��R�(KK��h�C
  �     �t�bhhK ��h��R�(KK	��h�C$p         M  	      	         �t�bhhK ��h��R�(KK��h�C       z   ,      X        �t�bhhK ��h��R�(KK��h�Cx     �  �   O     ;     I   %   /      �           �  �        �  C      �  h      �   �         �t�bhhK ��h��R�(KK��h�C\   w   �   �
              �     �       �        P      n      +         �t�bhhK ��h��R�(KK��h�CT
        2   �   0  p  
   z  �   7      �  �  p  
   z  s   7         �t�bhhK ��h��R�(KK��h�C1   #       �        �t�be.