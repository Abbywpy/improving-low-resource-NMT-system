Även i vår värld finns floder och träd och lejon och elefanter.
Står upp, går till ett hörn, den skälver,
Historien jag har berättat för er är stökig och oavslutad.
Central Intelligence Agency.
Låt oss leva med varandra och ta ett andetag i taget.
Det är en gentleman på första raden som faktiskt gör en exakt imitation av hur hon såg ut.
Vi vinner mark och snart kommer vi att övervinna krisen.
Hos de här barnen ville jag föra tanken till något som existerar inombords som ingen kan ta bort, så jag utarbetade en kursplan som dels är statsvetenskap, dels fotbollsturnering, i en konstfestival.
Det beklagliga är att våra städer, som New Delhi och Mumbai, inte har tillgång till vatten dygnet runt.
Ni kan om ni vill jämföra detta med, å ena sidan en hjärtinfarkt där man har död vävnad i hjärtat, kontra arytmi, där ett organ helt enkelt inte fungerar på grund av kommunikationsproblem inuti det.
Om du är ogift, sjunker siffran till tre.
Så detta är vad vi kallar en oktaeder.
Innan jag går vidare vill jag förtydliga min egen roll i detta.
Vi tog en annan grupp, en stor grupp amerikaner, och ställde en fråga i okunnighetens slöja.
Men, jag vet själv också, jag känner den här virtuella esprit de corps, om ni så vill, med dem allihop.
Vad pågår i den här bebisens huvud?
Kaffe både orsakar och motverkar cancer.
Den uppenbara frågan är, behöver verkligen ett TEDTalk 2300 ord?
(Applåder) CA: Under tiden, med hjälp av internet och den här tekniken, är du här, tillbaka i Nordamerika, inte riktigt USA, men Kanada, på det här sättet.
Verkligen inte. Låt oss se till att de närmsta 100 åren blir det bästa av århundraden.
Nummer 5: Osäkerhetsmomentet.
Jag skrev den här efter en väns begravning men inte så mycket om vännen som om något griftetalaren pratade om som alla griftetalare brukar göra, vilket är hur glad den avlidne skulle varit om hen tittade ner och såg oss alla samlade.
Doktor King trodde på att de fanns två typer av lagar i denna värld, de som skapas av en högre makt och de som skapas av människor.
Du ska till sydamerika, inte sant?"
(Skratt) Om jag går för långt åt andra hållet och gör det väldigt abstrakt vet ingen vad det är de ser.
Det här kanske ligger på gränsen till science fiction, men om även en liten del av det här scenariot blir sanning kommer vår ekologi och till och med vår art inte att klara sig länge oskadda ifrån det.
Så allt jag stoppade i min kropp ansåg jag vara medicin.
Ett av testen vi använde för kreativitet var alternativa användningsområden.
Jag arbetar med morgondagens forskare och ledare, och de förtjänar att få reda på vad vetenskapen säger så att de kan hjälpa till att forma en framtid för alla.
Beteendeekonomen Georg Lowenstein bad studenter på sitt universitet föreställa sig att få en passionerad kyss från en berömd person, vilken som helst.
Den var beviset på att jag inte hade räckt till, att jag var gammal och inte fantastisk och inte perfekt och inte passade in i den förutbestämda mallen.
Jag vet inget annat om honom, utom att han en gång räddade mitt liv genom att riskera sitt eget.
Vi behöver kunna säga någonting, för vet ni vilka fler som sitter vid bordet?
Han lyckades få till ett möte med fader Samaan, och överraskande nog älskade han idén.
Du ser att de som väntar till sista minuten har så fullt upp med annat att de inte har några nya idéer.
Men det provades aldrig.
Kära föräldrar, om ni skäms för mens, så kommer era döttrar göra det också.
Svar: Det tog dem, i genomsnitt, tre och en halv minut längre tid.
Och det är endast när vi hedrar dem och uppmärksammar dem och ger dem status som världen verkligen kommer att förändras.
Jag kom bara på besök och sade, "Det ser bra ut, bra jobbat," Det var allt. Ni kan se vad klockan är i alla fem kommuner av New York där bak. Så det här är utrymmet för handledningstimmarna.
(Skratt) Och en man kom att ge berättelser om sin far genom en plattform som heter Twitter för att kommunicera den skit hans far kom att uttrycka.
Det var en ordentlig utmaning, och det var faktiskt exempel från biologi som bidrog oss med många av ledtrådarna.
Varför vi väljer de semestrar vi väljer är ett problem vi möter med ett val mellan de två själven.
Och farmor, var fanns du när de marscherade med våra japansk-amerikanska grannar till interneringslägren?
Så låg inkomst här och hög inkomst här.
På andra områden snöar det eller så ökar ismassan igen på vintern.
Och om människor flyttar till urbana, okända, betongmiljöer så kan de också bli hjälpta i förväg av socialt stöd som redan väntar genom SMS-kunskap.
Trots det, 70 år senare, har cirkeln slutits.
Och i denna stund är vi perfekta, vi är hela och vi är vackra.
Bryr vi oss om människorna, vår familj, hälsa, eller är det prestation, framgång, sådant?
Sömnkvaliteten som du får som nattskiftsarbetare är normalt sett mycket dålig, återigen i femtimmarsregionen.
Det betyder inte att vi nödvändigtvis kommer till samma slutsats.
Han hade en mycket generös returpolicy, detaljerade köpvillkor, och kort leveranstid.
Och nu ska vi tända på det.
En dollar, tio dollar eller 100 dollar per dag.
Så snart den tilliten var uppbyggd ville alla vara med på vårt maraton för att visa världen Libanons sanna färger och det Libanesiska folket och deras önskan att leva i fred och harmoni.
Små finjusteringar kan leda till stora förändringar.
Så jag hoppas ni gillar det.
Det använder inte optik som ett vanligt mikroskop för att göra små objekt större. Istället använder den en videokamera och bildbehandling för att avslöja de minsta rörelserna och färgförändringarna hos saker och människor förändringar som är omöjliga för oss att se med blotta ögat,
Nu ser vi en stark ökning av nya konflikter och de gamla konflikterna är kvar: Afganistan, Somalia, Demokratiska republiken Kongo.
Jag var så hänförd av resultatet att jag ville plantera dessa skogar på samma sätt som vi tillverkar bilar, skriver programvara, eller driver vanliga verksamheter, så jag grundade ett företag, en end-to-end tjänst, för att skapa dessa inhemska naturskogar.
med den här inställningen. Den andra aspekten av min livsfilosofi är att jag omger mig med människor som jag vill vara med, människor av god kvalitet.
Vad alla dessa människor har gemensamt är att de är kättare.
Lunginflammation tog tre barn av tio.
Ta till exempel Airbnbs massiva succé som alla känner till.
I intervjun pratar hon med sin dotter Lesley om att som ung man gå med i ett gäng, och senare i livet bli den kvinna hon alltid var ämnad att bli.
För 150 år sedan beskrev anatomer väldigt, väldigt noggrant -- här har ni en modell av magväggen.
När en fluga rör sig över mittpunkten i kammaren där de två strömmarna av luktämnen möts, måste den ta ett beslut.
Och ingen skulle ge sitt livs besparingar till ökända smugglare om det fanns en laglig väg för migration.
Utförandezonen maximerar våra omedelbara resultat, och inlärningszonen vår utveckling och framtida prestation.
Och en sak man ser är att på manslinjen går dödligheten neråt, neråt, neråt, neråt, neråt.
Det var frihet under ansvar.
Innan vaccinerna fanns dödade många av infektionssjukdomarna miljontals människor per år.
Och det är mycket mer på gång.
Hon ville skapa ett bättre liv för sina barn och sin familj.
Om du verkligen bryr dig om att starta en rörelse, ha modet att följa och att visa andra hur man följer.
De är också silikon.
Jag är här för att berätta för er om framgång i Afrika.
Men finns det tänkbara händelser som kan vara ännu värre, som kan släcka ut allt liv?
Hur många av er använder skrivbordsfältet?
Undersökningsrummet kändes som ett skämt.
PM: Det tror jag inte. NA: Men det hjälper att berätta att några människor är agenter för förändring i samhället.
Som den där spindeln som bor bakom din soffa?
Men det är fortfarande lite komplicerat och lite svårt.
Mitt företag har mjukvara som gör detta redan idag.
Tack så mycket, Chris.
Jag undrade om vi kunde använda all data och all vår expertkunskap när vi utvecklar nätverk för att kvantifiera hur detta kan ske.
Men okej är aldrig okej.
För att nummer ett, svaret spelar roll.
Varje land i världen har tidningar. Den har ett bisarrt på pågående filosofisk projekt,
Så människor går omkring med virus som inte märks.
Dessa barn växer upp utan familjeförebilder eller en bild av goda föräldrar, så de kan ha svårt att själva vara föräldrar åt sina egna barn.
Detta är en plats av stor historisk betydelse.
Och om du drar på den här sidan av repet, försvinner repet från den andra sidan.
Vi ska inte oroa oss för vad våra maskiner kan göra idag.
Vi åkte tillbaka för den sista visningen av gården, och han visade mig de vilda pepparplantorna och växterna som han såg till fanns där för sältan.
Vår framtid är många-till-många.
Nyfikenhet och förundran, för den driver oss att utforska, för vi är omgivna av saker som vi inte kan se.
Det finns ingen som inte har gjort det så här långt.
Det är de blå staplarna.
Det var för fem år sen som jag verkligen började bryta ny mark genom att kombinera virtual reality och journalistik.
Så häng med mig runt och tillbaka i resonemanget.
Och det ledde sedan till mina stora frågor.
Ammoniaken avdunstar och den återkondenserar på andra sidan.
Just nu kan datorer göra det som människor ägnar det mesta av sin tid åt att göra för att få betalt, så det är hög tid att börja tänka på hur vi ska anpassa våra sociala och ekonomiska strukturer för att klara av den nya verkligheten.
Trots det är dessa miljöer bra platser för att stoppa den rörliga sanden.
Det förändrar hur du hanterar din upplevelse, det förändrar hur du tänker på din förövare, det betyder att om du träder fram, backar du upp någon annan och de backar upp dig.
Så livet måste förändras.
Så jag sprang ut i vinterkylan och fotograferade varenda person jag kunde få tag på i februari för två år sedan.
Lokal jihad blir global jihad igen om man struntar i det.
Hur löser då hjärnan sitt avfallsproblem?
Han fick sin arm amputerad för 10 år sedan.
Och vi beslöt att vi på minsta möjliga tid skulle förstå hur det nya viruset betedde sig i våra barn.
(Maskinröst) 1,8. Vi har många försök igång ute i byarna och i skolorna, och utifrån vad vi lärt oss ute i fält, har vi insett att det är viktigt att använda icke-medicinska termer så att människor kan förstå vad vi undersöker och vad det betyder för dem.
Och det verkar vara ett tryggt levnadssätt.
Så, på grund av den här explosionen i ljudtillgänglighet särskilt hos döva har detta inte bara påverkat hur musikinstitutioner och dövskolor behandlar ljud - och inte bara som terapimetod - fast som medgestaltare av musik, stämmer detta absolut också. Men det har betytt att akustiker verkligen har behövt fundera över vilka slags lokaler de konstruerar.
Flera år efter denna händelse tränade han racketbolltränarna.
För jag är kvinna.
Men en fantastisk person var han, en underbar filosof.
Det är en av de saker jag är mest stolt över i mitt liv.
Publiken: 23
Så jag säger till honom, helt klart i mitt huvud: "Det är Jill, jag behöver hjälp!"
När vi letar upp dem och frågar vad det är så säger de oftast något i stil med: "Jag är helt enkelt inte någon kreativ person."
Och när hon växte upp, när hon var fyra och ett halvt år gammal, skrev jag in henne i min skola.
En tid efter att den kom ut, väntade Augusten på en flygplats och besökte bokhandeln och tittade på vilka som köpte hans böcker.
Jag började med det för 15 år sen.
Och sen kom killen på en briljant idé, han sa, "Du driver ju den där organisationen Ungdomar Utan Gränser, eller hur?
Så jag tog reda på vad ekonomin betalade för kriget i Irak samma år.
Som många andra lägger jag mycket tid på att klaga över hur svårt det är att få människor att förändras, och vi borde inte tjafsa om det.
För när det gäller sex, är män pressade till att skryta och överdriva, medan kvinnor är pressade till att dölja, förminska och förneka, vilket inte är konstigt när man tänker på att det fortfarande finns nio länder där kvinnor kan avrättas för att de vänsterprasslar.
Förra året lyckades vi dock skrapa ihop lite pengar.
(Skratt) (Applåder) När vinden blåser, leds all överskottsenergi från vindkraftverket om till batteriet.
Att återta våra berättelser och lyssna på varandras, kan skapa en portal som kan överträffa tiden självt.
Som tur är så har vi en ny maskin, magnetencefalografi, som låter oss göra detta.
Uppmärksamhet är valutan.
Vi ser ett tydligt behov av att aktivt främja hälsoinsatser, särskilt bland äldre.
Jag har funderat och vägt samman hur det är att arbeta under kapitalism.
När han gör så, betyder det inte "Ta din Stradivarius och som Jimi Hendrix, slå den mot golvet."
Kometen är alltså fräsch och ny.
Det finns andra som nästan faller ihop när de kommer in, man ser det.
Var var den här för 10 år sen?
Folk vill alltid berätta saker om sina fantastiska skor.
Ändå spenderar vi överraskande lite tid för att ta hand om det som betyder mest: sättet vårt medvetande fungerar. Vilket, återigen, är det avgörande som avgör kvalitén på vad vi upplever.
När vi lär känna någon, lär vi oss hur de fungerar, och sedan lär vi oss vilka ämnen vi kan prata om.
Då kan vi börja använda celler.
Flickorna själva såg aldrig bilderna, men de gav dem till oss. Det är detta som kritikerna inte känner till, och det är denna forskning jag rekommenderar för de som vill arbeta humanistiskt.
Hon skulle antagligen säga att hon inte är så speciell, men hon har ett märkvärdigt inflytande.
Och, till skillnad från en massa choklad, kan massor av leenden faktisk göra dig friskare.
Det var inte okunnighet.
Jag var klar med skolan och skulle arbeta som juridiskt ombud och representera stammar runtom i landet, representera på Capitol Hill, och jag såg direkt varför rasistiskt bildspråk spelar roll.
Imorgon kommer det inte finnas någon ursäkt för att inte göra det rätta.
Och jag säger er att detta inte är en fråga om klimatpolitik eller miljöpolitik.
Och jag tänkte, jag ger dem ett prov. De kommer att få en nolla. Sen ger jag dem materialet. Jag kommer tillbaka och testar dem. De får en till nolla. Och går tillbaka tillbaka och säger, "Ja, vi behöver lärare för vissa saker."
Så fort som vi - och detta var på 50-talet - och så fort som vi tog bort det jagande, trummslagande folket för att skydda djuren, så började marken att försämras, som ni ser i den här parken vi skapade.
Så vi började prata om det här.
Detsamma är sant för genomskinliga solceller som är integrerade med fönster, solceller integrerade med gatumöbler, eller solceller integrerade med dessa miljarder apparater som bildar Sakernas Internet.
Till vänster har vi Casablanca, till höger har vi Chicago.
Om vi äter otillagad mat kan vi inte frigöra energin ordentligt.
Kort sagt spelar jag in en sekund av mitt liv varje dag i resten av mitt liv, och sedan i tidsordning sätta ihop alla dessa pyttesmå en-sekundare av mitt liv till en lång video tills jag liksom inte kan spela in längre.
Jag svarar, "Var inte oroliga, era föräldrar kan inte heller.
Ni känner alla till den här historien.
När män säger det handlar det ofta om något som de inte skulle ha gjort ändå.
Man filmar vägskyltar, klockor, dagstidningar.
Låt oss till exempel anta att det första fallet inträffar i Sydasien.
Det är inget fel på din hjärna. Det är inget fel på ditt förstånd. Du har Charles Bonnet-syndrom"
Revolutionen inom dödsvård har börjat.
Istället för att säga att det handlar om att vinna tävlingen, kommer folk inse att framgång mer handlar om att bidra.
Och uppfinningsrikedomen, om du nu kan kalla det för det, går djupare än så.
Det ligger på 826 Valencia Street i Mission-området i San Francisco, och när jag jobbade där låg högkvarteret för ett bokförlag där, som hette McSweeney's; en ideell skrivverkstad som hette 826 Valencia. Längst fram i huset låg en märklig affär.
Den använder de senaste molekylärbiologiska rönen, och är en billig, 3D-printad enhet, och datavetenskap för att försöka tackla en av mänsklighetens svåraste utmaningar.
Och hon bara: – Haha, något sådant finns inte.
I filmen "Spirited away" råkar de som tar emot guld från No-Face ut för otur.
Hon väntade otåligt på att flytta hemifrån. för att bevisa för dem att hon är vuxen, och för att bevisa för sina nya vänner att hon är en av dem.
Barnäktenskapen kommer kanske inte att bli färre.
Han är någon som flydde från allt detta dåliga."
Det är ett ställe vi går till för att komma bort från stressen i arbetslivet och ibland i familjelivet.
På franska till exempel skulle man säga "tu" när man pratar med sin kompis i skolan men "vous" när man pratar med sin lärare.
Det ni alla gör just nu med er bröstkorg, och sluta inte göra det, är att andas. Man använder interkostalmusklerna, musklerna mellan revbenen
Och deras kunder och miljön.
Vi följer dem som leder, inte för deras skull, men för oss vår egen skull.
Arkitekturens välbeprövade och genomtänkta formler och termer fungerar inte här.
Som resultat, tycker jag att vi stackars förtryckta kvinnor faktiskt har några nyttiga, surt förvärvade lärdomar att lära ut, lärdomar som kan visa sig användbara för den som vill blomstra i den moderna världen.
IndiGenomics handlar om vetenskap för folket och av folket.
Jag blev kallad en idiot, en förrädare, ett plågoris, en fitta och en ful man, och det var i ett och samma mail.
Man behöver inte en doktorsgrad för att se att det lämnar kvar 4 procent för resten av mångfalden.
Japan är världens äldsta land vad gäller snittålder.
Det stör mig eftersom jag varit öppen med min homosexualitet ganska länge nu.
Och för ett par år sedan bestämde jag mig för att skriva om prokrastinering.
Han bestämde att meningen med hans upplevelse var att få känna glädjen i vänskap och sedan lära sig att få vänner.
Och jag släpptes.
Hurra! Ni är grymma!
Jag hade ett konsultjobb tillsammans med en kollega och vi är så olika som två människor kan vara.
Och under nästa decennium kommer vi att ha ytterligare en miljard spelare som är extremt bra på vad det nu än är.
Det kan bli otroligt farligt när historier skrivs om eller ignoreras, för när vi förnekas vår identitet blir vi osynliga.
Deras konkurrenter är lika kvalificerade att göra alla dessa produkter.
Okej då, vad tror vi om det?
Vattnet blev hela min värld, varje krusning, virvel, näckrosblad och ström,
Tittar du för mycket på X Factor så köper du kanske idén om att alla kan bli vadhelst de än vill bli.
Jag vet inte hur Wagner lyckades med det.
Det kan du inte förvänta dig."
En av 20 personer röstade på vår kandidat som borgmästare i London.
Sperma som finns i kroppen i en vecka eller längre börjar utveckla avvikelser som gör att de inte är lika effektiva på att headbanga sig in i ägget.
Vi går tredje året på high school nu, och vi är mentorer åt yngre kårmedlemmar, som en enda sammanhållen grupp.
Detta är från Seattle.
Vi kan lära oss genom att iaktta andra människor och kopiera eller imitera vad de kan göra.
av respekt för de som kom innan en. Gå så här, tala så där, på grund av det.
Jag har skrivit en hel bok om det. Så jag lever för att lyssna.
Mumier är en fantastisk källa till information, men tyvärr är de geografiskt begränsade och begränsade i historisk tid också.
Varför inte ha den snabbtänkthet som Ken Jennings har, särskilt om man kan öka den med hjälp av nästa generations Watson-maskin?
Var så goda och delta i en tyst minut med mig.
Jag var orolig för dig när du sa att jag aldrig skulle lämna en tändsticksask någonstans i huset för att mössen kunde komma åt dem och starta en eld.
(Musik) Med era 2000-talsöron föredrar ni det sista ackordet, men förr i tiden skulle ni ha varit förbryllade, irriterade, och några av er skulle ha flytt rummet.
Men speciellt i USA väljer många unga bort att skaffa barn och det av samma anledning: ekonomisk oro.
Jag samlade pengar i Australien och återvände nästa år för att frivilligjobba på barnhemmet i några månader.
Och jag tror att det är högst osannolikt att de var långt från amerikanernas minne när de gick för att rösta i november 2008.
Det var en lögn, men det var min verklighet, precis som de bakåtsimmande fiskarna i lilla Dorothys sinne.
Men vi envisas med att förväxla objektivitet och subjektivitet som egenskaper hos verkligheten och objektivitet och subjektivitet som egenskaper hos påståenden.
De lärde oss hur man ger mediciner till möss.
Först gick det riktigt bra.
Svaret är, givetvis, att om man spenderar 125 miljarder eller 130 miljarder dollar per år i ett land, bjuder man in nästan alla,
Men underliggande makt är inte alls makt.
Och oavsett kultur, oavsett utbildning eller annat, verkar de här sju faktorerna vara närvarande när en person är i flow.
Jag är fortfarande exalterad över tekniken men jag tror, och jag är här för att lägga fram min teori att vi låter tekniken ta oss i en riktning, som vi egentligen inte vill.
Och det är bara fallet lån.
Och jag då?
Och den har utvecklats under tiden.
Ska vi vara oroliga?
Och på Stanford har man gjort sådan forskning i fem år nu för att dokumentera hur spelande med en idealiserad avatar förändrar hur vi tänker och agerar i verkliga livet, hur det gör oss modigare, ambitiösare och mer målinriktade.
Naturligtvis nyfikenheten, vetenskapsdelen av det. Det var allting. Det var äventyr, det var nyfikenhet. Det var fantasi.
Och ja, vi behöver hopp, det är klart vi gör.
Är de inte starkare?
och 100 företag utanför Idealab och försökte att komma fram till något vetenskapligt.
Jag överlevde på endast vatten.
Vi samlar blod från dem.
De är några av de minsta satelliter som någonsin avfyrats från världens största satellit.
Hur förändrar vi transportvägarna - för varor och människor?
Vi har två väldigt tävlingsinriktade, datakunniga företag.
Det är en invecklad dans i 28 000 km/h mellan vår kapsel, som är lik en pytteliten bil, och rymdstationen, som är stor som en fotbollsplan.
Många av oss går genom livet och försöker göra vårt bästa i allt vi gör oavsett om det gäller arbetet, familjen, skolan eller något annat.
(Applåder) Jag har utlovats förändring sedan jag var barn.
Det var mycket svårt, ska du veta, att göra min auktoritet gällande.
Om vi stabiliserar sömnen hos de individer som ligger i riskzonen så kan vi helt säkert göra dem friskare men också lindra vissa av de förskräckliga symptomen hos mentala sjukdomar.
För ur den urbana förstörelsen i Port-au-Prince kom en storm av SMS, människors rop på hjälp, bönfallandes för vårt stöd, delandes information, erbjudandes hjälp, letandes efter deras nära och kära.
Var jag än kom, kände det som att min fantasi, var den enda resväska jag kunde ta med mig.
Deras biblar har en liten inskription, det står "USA:s armé" på dem.
Och jag antar att du injicerar det kanske i ett strutsägg, eller något sådant. Och sedan väntar du och, hör och häpna, ut poppar en liten dinosaurieunge.
Gatorna översvämmades men folk ville inte missa chansen att delta vid en sådan nationaldag.
(Skratt) Varför framhärdar vi med att göra samma sak om igen och ändå förvänta oss olika resultat?
Briljant!
När uppgifterna kom tillbaka räknade jag ut betyg.
När detta gjordes - jag ber om ursäkt - jag kommer använda en förlegad jämförelse mellan uppslagsverk och Wikipedia, men jag gör det för att peka på att när vi gjorde denna inventering, var vi tvungna att titta på massiva mängder information.
Och i allra första början är inte alls så många berörda. och då får den klassiska sigmodala, eller S-formade, kurvan.
Så det är detta som används.
Så att fly från det verkliga samtalet kan ha betydelse eftersom det äventyrar vår förmåga till reflektion.
En tredjedel av alla frukter som vi äter är ett resultat av att insekter tar hand om växternas reproduktion.
De kommer behövas för arbete med avancerade skattefrågor och avgörande stämningar.
Men det finns en art i Everglades som du, vem du än är, inte kan låta bli att älska, och det är rosenskedstorken.
Varje dag bygger alla vi här gudar som har blivit alldeles vildvuxna, och det är dags att vi börjar slå ner dem och glömma deras namn.
Väck dina åhörares nyfikenhet.
Under en lång tid har människor sett vetenskap och humaniora som åtskilda.
Vilket jag tycker var en intressant idé, teori.
Och detta, så klart, är grundvalen i mycket av den österländska filosofin. samt att det inte finns något oberoende Själv, skild från andra mänskliga varelser, som inspekterar världen, inspekterar andra människor.
Tio år senare, en annan historia: Iranska revolutionen 1979.
Nuförtiden får ett av 88 barn diagnosen autism, och frågan är varför kurvan ser ut på detta sätt?
Vi gör detta genom att tänka igenom veckan innan vi befinner oss i den.
Där, mina damer och herrar, utvecklas den amerikanska demokratin under Thomas Jeffersons hand.
Okej, så vad är synestesi?
(Skratt) Desto smalare jag blev, desto längre kunde jag hålla andan.
Om civilbefolkningen dödas, om vapnen tar sikte på samhällen kommer det att föda en ond cirkel av krig, konflikt, trauma och radikalisering och den onda cirkeln är mittpunkten av så många säkerhetsutmaningar som vi står inför idag.
(Skatt) Så för att ta tag i problemet samlade jag en grupp internationella forskare i Schweiz, Danmark och Storbritannien
Idag tycker jag datorer gör motsatsen.
Jag skapar bilderna genom att välja bland korten i ett massivt arkiv från satellitföretaget Digital Globe.
Håll upp den.
Jag har identifierat mig på olika sätt - som bisexuell, som lesbisk - men för mig innefattar queer alla lager av den jag är och hur jag har älskat.
Vi var ense om att adresser är dåliga.
Min etik för att iaktta är formad av 25 års erfarenhet av att rapportera om tillväxtekonomier och internationella relationer.
Och när jag säger "väldigt vanligt" kan det fortfarande vara så sällsynt att inte en enda ö av liv någonsin möter en annan, vilket är en sorglig tanke.
Så den kvällen, la jag ut det på Facebook och frågade några av dem, och på morgonen hade svaret varit så överväldigande och positivt, att jag visste att jag måste prova.
Syntetisk biologi, till exempel, strävar efter att beskriva biologi som ett designproblem.
Vi måste omdefiniera i grunden vilka som är experter.
Hon var dotter till människor som faktiskt varit slavar.
Det hade pH 11, och ändå levde kemosyntetiska bakterier i det. I denna extrema miljö.
Vi är inte färdiga med videon än.
När du rör din arm så här, skickar hjärnan en signal till dina muskler här.
så tänker jag "nej, nej, jag vill inte ta konstgjorda preparat, jag vill bara se växter och - bara visa mig örter och växter. Jag vill se alla naturliga ingridienser".
Vissa är mindre.
Men duvan, som uppenbarligen aldrig gick i flygskolan, sprattlar till, flop, flop, och landar på ena änden av min balansstång.
Det är under sömnen vi återställs och återuppbygger oss själva, och när ett hotfullt buller som det här håller på, säger din kropp, även om du lyckas somna, så säger din kropp till dig: "Något hotar mig. Det här är farligt."
Föremålet som formade detta var troligen mellan 30 och 50 meter tvärsöver, vilket grovt sett är storleken på Mackeyauditoriet här.
vilket betyder att du kan skapa mening och bygga identitet och fortfarande vara fullständigt ursinnig.
Ni? OK. Först av allt, vilket år var det?
200 miljarder baspar i veckan.
Psykoanalytisk psykoterapi fyra-fem dagar i veckan i decennier och fortlöpande, samt utmärkt psykofarmaka.
Ett svar min fru kunde ha gett.
Rättigheterna vinns inte i rättssalar, utan i människors hjärtan och själar.
Det skulle bli ett köpcenter, istället för en grön oas.
Vi kallar varje avläsning för en emotionell datapunkt, och de kan aktiveras tillsammans för att visa olika känslor.
Men en sak jag är riktigt nervös för är mina skakande händer.
Jag växte upp med en mycket berömd farfar, och vi hade en sorts ritual därhemma.
LED-lampan strömmar nu videon genom att ändra dess ljusstyrka på ett subtilt sätt. ett sätt som inte uppfattas med vanlig syn, eftersom förändringarna sker för snabbt för att märkas.
Det här slog mig när jag skulle köpa nya jeans.
I Ryssland anses jag vara en gammal nucka som aldrig kommer att bli gift.
Och att man inte kan existera i det här universumet utan massa.
Ritualerna var bekanta.
Och jag tror att TV:n är som en global lägereld.
I kvantvärlden behöver du inte kasta den över muren, du kan kasta den mot muren, och det finns en viss icke-noll sannolikhet att den försvinner på din sida och dyker upp på den andra.
Ta, till exempel, ljudet av ett skott.
Vi kommer inte att bryta med dig, och det är något jag alltid har velat att du ska veta, att du är älskad.
Det har gett oss motivation till att fortsätta att jobba på detta.
Så bara en vecka efter Bergenbanan, ringde vi företaget Hurtigruten och började planera för nästa program.
Jag är inte en religiös eller särskilt andlig person, men i vildmarken, tror jag att jag upplevt religionens födelseplats.
(Skratt) Inte för att jag är en dålig lärare, utan för att jag har studerat mänskligt avfall och undervisat i hur avfall transporteras genom reningsverk, och hur vi bygger och designar dessa reningsverk för att skydda ytvatten, till exempel floder.
Det var en rätt fantastisk upplevelse, men det är fyra år sedan nu.
När du kombinerar vetenskapen bakom att känna igen bedrägeri men konsten att titta, lyssna, befriar du dig dig från att samarbeta i en lögn.
SM: Ah, ett drag av klassisk övervakningsekonomi.
Han bodde i ett område med få vägar där det rådde en stor brist på sjukvårdare.
Extas är alltså att man går in i en alternativ verklighet.
Vi kyler ner våra system till nära absoluta nollpunkten, vi utför våra experiment i vaakum, vi försöker isolera dem från alla yttre störningar.
Men har vi nått vårt mål?
Vi kan surfa på nätet anonymt.
I stället var det min välsignelse och förbannelse att bokstavligen bli människan i tävlingen mellan människa och maskin som alla fortfarande pratar om.
När vi funderar över konsekvenserna av det och vi tror på att utrotning är vanligt och naturligt normalt och uppstår då och då blir det i högsta grad moraliskt rätt att ha en mänsklig mångfald.
Så jag ber er att sprida informationen och håll ögonen öppna.
Ett ärligt svar för några månader sedan hade varit, "Vi har ingen aning."
Thailand, 64 procent.
På Comic-Con eller någon annan Con fotar man inte bara folk som går omkring.
Men sedan förstod jag, det är det redan.
Lycka till den här veckan.
Jag skulle vilja lägga denna typ av fredagskväll-i-baren-diskussion åt sidan och få dig att faktiskt kliva in i labbet.
Fienden har en röst.
Gör som jag, är ni snälla.
2004 så producerade de amerikanska drönarna totalt 71 timmar övervakningsvideo för analys.
Studenterna åkte dit i förväg, och de ordnade så att alla skulle beställa Feynman-smörgåsar.
Och dagar har blivit till månader, månader till år.
Jag fick lämna dem utan ett ordentligt avsked.
"Oh förlåt, jag blev lite sen. Hur går det?"
Äktenskapsmäklaren tänkte igenom allt, sammanförde två personer, och så var det bra med det.
Jag säger "Gud, jag önskar verkligen att jag hade kopplat ihop John Locke's teori om äganderätt med de efterföljande filosoferna"
Om vad?
Och du borde ha alla nätverk från alla dessa relationer mellan dessa element av data.
Och nu har vi många bakteriestammar i vår frysbox som får koraller att gå genom den där bosättningsprocessen.
Vi reste till byn för att mobilisera samhället.
Min fru började bötfälla mig på en dollar för varje irrelevant fakta jag förde in i vår konversation.
Eleven försökte, lyckades nästan, men fick det inte att bli alldeles korrekt.
Och du har inte varit dig själv.
Landskapet har sorgligt nog befolkats med fler fall som mitt, oavsett om någon har gjort ett misstag eller inte, och nu berör det både offentliga personer och privatpersoner.
Att bli blind satte dem i fokus.
Ryan Holladay: Blanda utan skarvar.
Och det kanske låg lite sanning i det där, för jag trodde att om jag bara började gå så skulle alla andra, ni vet, följa med.
I filmer är det helt annorlunda.
(Skratt) Och sedan odlade vi celler på dem.
Du kan alltså ha inte bara "bilceller", utan "Aston Martinceller"
Mitt sätt behöver dem inte.
Människorna.
(Musik) God eftermiddag.
Men mycket viktigare, fördelningen är mycket bredare.
Redan som barn förstod jag vilka förväntningar som fanns på mig.
Jag var inte för juridik.
Den har allt inbyggt, och den hoppade för att en student tände en bordslampa bredvid den.
De kommer att vara tillgängliga via maskinen.
Datan visade att jakten på lycka kan göra människor olyckliga.
Så därför. Om du ser här, nu kan jag fortfarande se det.
De jämförde Dreyfus handstil med den på anteckningen och drog slutsatsen att de stämde överens, även om professionella handstilsexperter utanför det militära var mycket mindre övertygade om likheten, men strunt i det.
KKM: Jag har tvingats påminna mig om en massa saker, jag också.
Vi behöver tusentals åklagare för att se detta och skydda dem.
Men om vi kan få den data ut från bakom fördämningen så att mjukvarutvecklare kan hoppa på dem, på det sätt som dessa utvecklare gillar att göra, vem vet vad vi då kommer att få fram.
Mitt favoritexemple är en borrmaskin. Vilka här äger en borr, en hemmaborrmaskin?
Vi fick veta att han hade en lång bakgrund av våld i hemmet.
Missförstå mig inte, det vore jättehäftigt att hitta utomjordingar.
Här fattas just nu beslutet att du förmodligen inte kommer beställa stek till middagen.
Det är ett praktexempel på vad som händer när regeringar attackerar deras egna medborgare. DigiNotar är en certifikatutfärdare
Tyvärr är det inte slutet på historien.
(Skratt) CA: Sa han att du skulle hoppa, eller var det mer som "Jag drar nu!
de är faktiskt skadliga.
och du log mot den jävla kameran som de sa till dig att göra eller så kunde du kan säga hejdå till din födelsedagfest. Men ändå, jag har en enorm stapel
Det finns människor - några har jag redan nämnt - som är fantastiska, som tror på kvinnors rättigheter i Saudiarabien, som försöker och som får ta mycket hat eftersom dom tar ton och gör sig hörda.
Men det finns 22 länder där man talar arabiska och de använder modern standardarabiska, som är den arabiska som används i hela regionen i tidningar och i TV och radio, men självklart skiljer det sig åt mellan länderna i vardagsspråket i dialekter, vardagsuttryck, och så vidare.
Vi kan kalla honom Miguel. Hans namn är faktiskt Miguel.
(Jag är hungrig!)
De får dig att betala mer i källskatt bara för att bättra på deras pengaflöde.
Här är ett foto på mig - jag är överlycklig.
Icke-statliga organisationer förstår fördelarna med att ha reportar som följer deras arbete vid sidan om.
Trappistmunken Thomas Merton frågade under Apolloperioden, "Vad kan vi vinna på att segla till månen om vi inte förmår korsa avgrunden som skiljer oss från oss själva?"
Vi behöver transformerande förändring.
Den klimatrelaterade extrema torkan som började 2006 i Syrien ödelade 60 procent av jordbruken i Syrien, dödade 80 procent av all boskap, och tvingade 1,5 miljoner klimatflyktingar till Syriens städer, där de kolliderade med ytterligare 1,5 miljoner flyktingar från Irakkriget.
För att lyckas behöver vi alla tillsammans hjälpa och påverka våra politiker, eftersom utan långtgående, världsomspännande förändring så kommer det inte att hända något.
Istället säger de. 'Nej, nej nej!
I Bangladesh finns ett område som heter Matlab.
Året efter, 1949, gjorde vi beslutet permanent i den nya författningen, och det är därför jag kan berätta denna historia nästan 70 år senare.
(Skratt) Just nu har vi väldigt lovande pilotdata.
Vi använder förstås elektricitet. Men vi har en lösning åt er - Vi använder oss av en ren energikälla.
2000 år senare kan vi förklara vad som händer i hjärnan.
Om vi gör så här tillräckligt ofta, och vi gör det med respekt, kommer folk att tänka efter lite mer kring hur de sätter ihop mötesinbjudningar.
Jag frågade dem varför.
En gång tvittrade jag, var i Lembourne kan jag köpa en netiflaska?
Det här är Emma Ott.
Och vi kommer bara att bli tio miljarder i världen, om de fattigaste människorna kommer ur fattigdom, att deras barn överlever och att de får tillgång till familjeplanering.
Istället för att arbeta i samklang med min omgivning, motarbetade jag den.
En garderob är bara ett svårt samtal och även om våra ämnen varierar oerhört mycket, så är upplevelsen av att vara i, och komma ut ur garderoben, universell.
Det var en plåga.
Så tänk om jag istället för att låta folk summera enskilda TEDTalks till sex ord, gav dem 10 TEDTalks på en gång och sade, "Sammanfatta dessa med sex ord åt mig."
Snart, hoppas vi, ska Masa få återförenas med honom i Sverige, tills dess tas hon om hand på ett vackert barnhem i Aten.
Det är faktiskt så att antalet människor som är inblandade i att tillverka en bil har ändrats ytterst lite de senaste årtiondena, trots robotar och automation.
Donald gav oss några av dessa läxor.
Skulle vi använda vår auktoritet och makt för att försöka kontrollera eleverna för att hindra dem från att gå, eller skulle vi stötta dem då de utövade de principer om social rättvisa som vi undervisat om sedan årskurs 9?
Och en av dem är att jag klarar mig bra.
Men det är en enorm skillnad mellan Afghanistan och Sri Lanka.
Okej, så ni förstår tanken.
Kan det stämma? Det gör det. Han var 33, 38 och 63 när de gjordes.
Och den här tävlingsretoriken är standard nu.
Men man kan bygga ett godtyckligt antal tunnlar, hur många nivåer som helst.
Och sedan byggde hon huset.
För jag vet inte om det finns något värre när det gäller den globala folkhälsan än att låta barn på denna planet dö av sjukdomar som kan förebyggas med vaccin, vaccin som kostar en dollar.
Så vi vet att de här kråkorna är riktigt smarta, men ju mer jag grävde i det här, ju mer upptäckte jag att de har gjort en till och med ännu viktigare anpassning.
Låt mig gå igenom dessa tre saker.
Män drabbas av autism fyra gånger oftare än kvinnor och vi kan verkligen inte förstå vad som orsakar detta.
De tappade lusten långt innan de har kommit hit.
Jag minns att mina sköterskor klagade på att köra genom det.
Spejaren är den som går ut, kartlägger terrängen och identifierar potentiella hinder.
Varför designar jag inte något som mäter fuktnivån i såret så det kan hjälpa läkare och patienter att behandla såren bättre?
Även om vi kunde mäta vad varje cell gör i varje givet ögonblick, måste vi fortfarande få ordning på mönstret i den inspelade aktiviteten, och det är så svårt, risken är att vi kommer förstå precis lika lite av dessa mönster som hjärnan som producerar dem.
Vi ska göra detta på människor som har kognitiva störningar och vi valde att behandla patienter med Alzheimers som har kognitiva brister och minnesförlust.
De försvinner på grund av att vissa företag inom skogssektorn går in och skövlar allt.
Det var det vanligaste svaret som vi fick.
och istället för att använda magneter eller muskler för att få den att röra sig så använder vi raketer.
Leopardsälen har sedan Shackletons tid haft dåligt rykte.
När jag studerade i Italien, insåg jag att jag saknade arabiskan.
Och i en bakterie gör CRISPR-systemet det möjligt att plocka ut DNA:t från viruset och integrerat i små bitar in i kromosomen - i bakteriens DNA.
Den ena är att de är mycket vanliga.
Så två saker i det här slog djup an hos mig.
Nummer ett: Vi måste börja göra våldsbekämpningen till en självklarhet i kampen mot fattigdom.
Och deras ledare, deras ledare: innan de skickar sina söner och döttrar att kriga i ert land - och ni vet varför - innan de skickar iväg dem går de till en kristen kyrka och ber till sin kristna gud och ber om skydd och vägledning från den guden.
De föddes alla in i den eller så har de aktivt strävat efter att omge sig med rätt folk.
Så medlemmar i mitt team reste omedelbart ut och anslöt till Dr. Humarr Kahn och hans team, och vi möjliggjorde för diagnostisering med känsliga molekylära tester för att fånga upp ebola vid gränsen in till Sierra Leone.
Att acceptera det faktum att vi är djur får en del potentiellt skrämmande konsekvenser.
Om man tar någon som Portia de Rossi, till exempel, så är alla överens om att Portia de Rossi är en mycket vacker kvinna.
Räck upp en hand om du är i 20-årsåldern.
Det var så, kreativiteten måste hitta sitt utlopp på något sätt.
Ute i världsrymden har vi nu en människotillverkad sattelit, som uppenbarligen sänder ut någon slags signal. Om vi hittar rätt våglängd kan vi nog höra den."
Jag började ta fram en ny typ av fjärrstyrning. Med robotars hjälp kunde jag vara på flera ställen samtidigt- -utan att behöva ta mig dit själv.
Notera bokens titel, "Boken som aldrig checkades ut: Titanic."
(skratt) Jag tänkte "Ja, det är fantastiskt, för jag känner mig inte handikappad".
jag blev tvungen att leva med två helt olika bilder av mig själv som person; som en skurk hemma i mitt hemland och som en hjältinna i världen utanför.
När Patrick kom ut från fängelset hade han en olidlig resa framför sig.
Jag har investerat i Pakistan i över sju år nu, och de av er som också arbetat där kan skriva under på att pakistanier är en otroligt hårt arbetande folk, och det finns ett häftigt avancemang uppåt i deras natur.
i vårt land. För ytterligare bevis kan vi se på fängelsestatistik; vi kan se på statistiken över polisvåld gentemot svarta; vi kan se på utbildningsklyftan - så ja, social rättvisa hör hemma i skolan.
30 färdigheter kunde rädda 30 miljoner liv före år 2030.
Krigets framtid innehåller också en ny typ av krigare, och det håller faktiskt på att omdana upplevelsen av att gå i krig.
Vi har än så länge inga genetiskt förändrade människor, men det är inte science fiction längre.
Som vanligt talade vi om världsproblemen.
Och mitt absoluta favoritord inom denna kategori är "multi-slacking".
Hon har faktiskt en Harvardpsykolog och har behandlats för bland annat affektiv sjukdom
Man behöver inte gå till apoteket längre.
Om vi nu vill undersöka detta närmare?
Det sista landet – det sista landet i världen som avskaffade slaveri är samma land som jag föddes i, Brasilien.
Varför kände jag mig så berättigad att döma henne?
Jag behöver vila den här veckan," eller "Jag behöver crossträna.
Alldeles strax kommer ni höra ett tåg som de inte reagerar på.
Det fanns inga incitament för någon att förbättra produkten, eftersom den finansierades av gåvor.
Och det är möjligen de största som någonsin hittats.
Så när jag tänker vad som är det fundamentala värdet av ett företag som Tesla, skulle jag säga, förhoppningsvis, om den påskyndade processen med ett decennium, möjligen mer än ett decennium skulle det vara en väldigt bra grej.
Så vi måste ställas inför denna fråga: hur får vi våra 1900-talslagar för krig, som är så åldersstigna nu att de har rätt till äldrevård, att hinna ikapp denna teknik från 2000-talet?
Vi vet till exempel, från forskning, vad som är viktigast för de som är nära döden: komfort; att känna lättnad, att inte vara en börda för sina kära; existentiell frid, och en känsla av förundran och andlighet.
Se bara på de här vackra, fascinerande varelserna.
Ni förstår vikten av det?
Och ni användare; det gäller oss alla - vi kan kräva teknik som fungerar på det här sättet.
Men, jag hoppas att ni håller med mig om att dessa saker som jag precis beskrivit för er, var och en av dem, förtjänar någon form av pris. (Skratt) Och det är vad de fick, alla fick ett Ig Nobelpris.
Brutus är Venus granne och "ställa till med bråk" är det som hände dagen efter Venus man hade dött, när Brutus bara kom och slängde ut Venus och hennes barn från huset, stal deras mark, och rånade deras marknadsstånd.
Mitt dysfunktionella själv kunde faktiskt koppla in till ett annan själv, inte mitt eget. Och det kändes så bra.
Med åren har verktyg blivit mer och mer specialiserade.
Där finns inga stora gravkammare som de flesta kyrkogårdar kräver bara för att formgivningen ska bli lättare för dem.
Jorden kan sedan användas till att skapa nytt liv.
Jag vet inte." Ni vet vad det innebär.
Dina minnen och associationer och så vidare.
(Skratt) Arton minuter, uppenbarligen omöjligt.
Den till höger är den som får vindruvor.
Du verkar tröttna Bob, men håll ut, för här är den verkliga superegenskapen.
Och om vi inte lägger tid och uppmärksamhet på det och tillgodogör oss det lärandet och applicerar det på resten av livet, då är det meningslöst.
Men de tävlar även efter att de parat sig, med sin sperma.
Detta visade sig vara mycket värdefullt 20 år senare då Michael Bloomberg bad mig bli hans stadsbyggnadschef och gav mig ansvaret att omforma hela staden New York.
Min "Svart kille"-grej är så bred och så djup att jag i princip kan sortera och lista ut vem den svarta killen är, och han var min svarta kille.
De är som biologiska fönster som lyser och berättar att cellen nyss var aktiv.
Allt började i vårt garage.
Här är hon, en Hollywoodkunglighet. Jag är en tuff unge från Detroit, [Dolly] är en sydstatsunge från en fattig stad i Tennessee, och vi fann att vi var så synkade som kvinnor, och vi måste ha - vi skrattade - vi måste ha lagt till åtminstone ett årtionde på våra liv.
Jag kunde rita. Jag kunde måla.
Och jag tror att när du söker efter ledarskap, måste du se inåt och mobilisera ditt eget samhälle för att skapa förhållanden som öppnar för en ny sorts lösning.
Den värms upp under cirka 30 minuter, kyler ned på ungefär en timme.
Dopaminet som strömmar runt när du är positiv, har två funktioner. Det gör dig inte bara lyckligare,
Dessa bilder från American Society for Microbiology visar oss processen.
Den första är floden av data som skapas av drönare.
Som någon som är ganska nära världsrekordet i antal timmar som tillbringats under en magnetkamera kan jag berätta att en förmåga som är väldigt viktig inom MRT-forskning är kontroll över blåsan.
Jag deltog i ett seminarium i år med en skådespelande lärare, Judith Weston.
Och det andra alternativet som kan bli klart i tid är hushålls-solel kompletterat med naturgas, vilket vi kan använda i dag, kontra batterierna som fortfarande är under utveckling.
"Har du nånsin träffat nån som vaknat på morgonen - (Skratt) och blivit svart?"
Tanken var -- med samma utgångpunkt, ett splittrat land -- att samla tecknare från alla läger och låta dem skapa något tillsammans.
Så det är bra, men naturligtvis skulle vi ännu hellre hitta ett sätt att påverka funktionen i hjärnregionen, och se om vi kan ändra på människors moraliska omdömen.
Detta var bakslaget i Kenya och Ghana gick förbi, men sedan dalar Kenya och Ghana tillsammans. Fortfarande stillestånd i Kongo.
Det finns fler: habitatförlust är en av sakerna jag ofta bryter ihop inför mitt i natten.
För mig är de pillren analogin till bilstolarna.
Hon säger att det inte finns något mer sinnligt än en het dusch, att varje vattendroppe är en välsignelse för sinnena.
