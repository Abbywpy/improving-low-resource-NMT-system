återbetalas (1/1)
industrin (1/1)
musikinstitut (3/3)
medium (1/1)
korttidsrehabilitering (1/1)
kortti (2/2)
nummerserie (1/1)
kommunerna (18/18)
utöva (8/8)
A2.2 (1/1)
dyrt (1/1)
kollaps (1/1)
potilasasiamies (2/2)
parentes (1/1)
sakkunniga (1/1)
patientens (2/2)
kansli (7/7)
kedja (1/1)
Vailla (1/1)
alternativa (1/1)
medborgarskapsanmälan (4/4)
bankernas (1/1)
precis (2/2)
studielån (4/4)
näringsbyrå (14/14)
anställning (21/21)
bostadsaktiebolaget (6/6)
gynekologisk (1/1)
läkarrecept (3/3)
työttömyyskorvaus (2/2)
material (13/13)
platser (5/5)
solen (3/3)
anmält (4/4)
kommunen (34/34)
föräldraskapet (4/4)
skolkuratorn (2/2)
pappersformulär (1/1)
försäkringar (9/9)
insamlingsställen (1/1)
Hyvin (1/1)
friluftsleder (1/1)
boendeform (1/1)
förete (1/1)
avfallet (5/5)
vidimerad (1/1)
yrkeskunskap (1/1)
Sportkort (1/1)
storfurstendömets (1/1)
starta (17/17)
sjunger (1/1)
förvärvats (1/1)
träsliperi (1/1)
aikuiskoulutustuki (1/1)
betalningskrav (1/1)
konkurrerar (2/2)
civilvigsel (1/1)
yrkesexamen (11/11)
registrerade (6/6)
telefonsamtal (1/1)
utevistelse (1/1)
hemsjukvården (1/1)
yhdessä (1/1)
avgiftningsvård (1/1)
bostadsrättskontraktet (1/1)
uppehålla (1/1)
sökfält (1/1)
redogörs (1/1)
trottoaren (1/1)
guiden (2/2)
tasa (2/3) Tasa (1)
perhe (1/1)
TTS (1/1)
kommunicera (1/1)
häva (2/2)
menas (1/1)
Åboregionen (1/1)
förändringar (2/2)
vise (1/1)
skaffa (26/26)
åldersspannet (1/1)
värmeelement (1/1)
hälsostationens (1/1)
besvärstillstånd (2/2)
löper (4/4)
Ajovarmas (2/2)
konstruktionen (1/1)
läroavtalsutbildning (5/5)
vigseltillfället (1/1)
organisationers (2/2)
mat (18/18)
läder- (1/1)
obetald (1/1)
vån (14/14)
människogrupp (1/1)
rundvandringarna (1/1)
vaccination (1/1)
personefterforskningen (1/1)
läkemedelsbutikerna (1/1)
peruskoulu (3/3)
frysens (1/1)
aikuiskoulutuskeskus (1/1)
inriktning (1/1)
formen (1/1)
pauserna (1/1)
fylla (19/19)
per (60/60)
hälsovårdstjänsterfinska (1/1)
kök (1/1)
centralt (1/1)
körning (1/1)
avslutade (2/2)
far (9/9)
hörde (2/2)
ylempi (1/1)
Ingående (2/3) ingående (1)
hengenvaara (1/1)
infödda (1/1)
tvättmaskinen (1/1)
yrkesskola (1/1)
stadshus (2/2)
yrkesutövning (2/2)
färdigheterna (1/1)
Rovaniemen (2/2)
krisjourenfinska (2/2)
vägledning (5/5)
möbler (4/4)
arbetspensionssystemet (1/1)
stor (10/10)
start (1/1)
euro (23/23)
handeln (4/4)
varför (4/4)
intervju (1/1)
fördela (2/2)
digitalbox (1/1)
reparationer (5/5)
nordiskt (7/7)
täckande (1/1)
vanligtvis (47/47)
kända (1/1)
kung (4/4)
full (4/4)
boningsort (1/1)
dig (368/368)
återflyttare (2/2)
straffa (1/1)
billigast (1/1)
sättet (4/4)
tullmyndigheterna (1/1)
chefen (1/1)
Inkomstregistrets (1/1)
Helsingforsfinska (9/9)
sjöar (1/1)
mångformigt (1/1)
ungdomspsykiatriska (1/1)
anställningsintervjun (1/1)
jordbruks- (1/1)
arbetssökning (1/1)
Tyskland (1/1)
föreskrivs (2/2)
parkgympa (1/1)
byta (8/8)
tämligen (1/1)
vuxna (33/33)
illegalt (1/1)
lastenneuvola (5/5)
researrangemangen (1/1)
nödsamtal (1/1)
samhälleliga (1/1)
uppsökande (3/3)
fientlig (1/1)
tillstånden (1/1)
presidentens (1/1)
dock (54/54)
dröjsmålsränta (1/1)
görs (37/37)
tillåter (3/3)
denna (22/23) Denna (1)
stadsbor (1/1)
överinspektören (1/1)
vägnar (1/1)
vederlagets (1/1)
hyresetta (1/1)
invandrarfamiljer (1/1)
påbyggnadsutbildning (4/4)
veckovisa (1/1)
responssystemet (1/1)
personligen (11/11)
bostadsrättsavgift (1/1)
jour (1/1)
rullstol (1/1)
Internetfinska (8/10) internetfinska (2)
Naiset (1/1)
anmäler (14/14)
politiska (6/6)
utredningen (3/3)
förlora (7/7)
ägo (1/1)
Pensionsskyddscentralens (1/1)
upprättas (5/5)
fort (8/8)
sju (8/8)
bodelning (1/1)
undervisningssektorn (1/1)
dödsorsaken (2/2)
oavlönad (3/3)
arbetsinkomsten (1/1)
innebär (20/20)
judiska (1/1)
psykisk (3/5) Psykisk (2)
asylansökningsblankett (1/1)
kurser (36/36)
utrikespolitik (1/1)
överenskomna (2/2)
medlemsländerna (1/1)
bostadsbidrag (20/25) Bostadsbidrag (5)
museets (1/1)
FRK:s (1/1)
Twitter (1/1)
skyddfinska (4/4)
papprullar (1/1)
espoo.fi (1/1)
klassificerats (1/1)
spelberoende (3/3)
arbetslöshetskassor (1/1)
budget (1/1)
mete (1/1)
Yrkenas (1/1)
eget (62/62)
systerdotter (1/1)
ersätta (8/8)
bilplatser (1/1)
pensionsinkomster (1/1)
olyckor (2/2)
studiestödfinska (1/1)
tron (2/2)
investerare (1/1)
UNHCR (4/4)
konstruktioner (2/2)
utställningar (7/7)
skäl (14/14)
beordra (1/1)
verkställa (1/1)
organisationens (2/2)
antal (4/4)
anser (3/3)
medicinskt (1/1)
studera (89/89)
byggbranschen (1/1)
klädregler (1/1)
damm (1/1)
tim. (1/1)
hemtjänster (1/1)
biometriska (1/1)
besvären (4/4)
skulder (10/10)
fukt (2/2)
rutt (4/4)
slutat (1/1)
hygienpass (1/1)
länge (27/27)
ökar (1/1)
erityisammattioppilaitos (1/1)
subventionerade (1/1)
finansiärer (2/2)
opetustoimi (1/1)
idrottsväsendet (1/1)
befunnit (1/1)
tillgängliga (3/3)
avlönat (1/1)
näring (1/1)
pris (6/6)
dagvårdplats (1/1)
ansvara (1/1)
smälter (1/1)
Suomenkielisen (1/1)
ville (2/2)
universitetfinska (6/6)
procent (26/26)
friluftsliv (4/4)
gjorda (1/1)
Tammerfors (2/2)
kommunala (18/18)
banklån (4/4)
jurister (4/4)
avtalad (2/2)
ute (3/3)
www.tuotos.fi (1/1)
bilagorna (4/4)
öppnas (1/1)
porten (1/1)
ungdomsgårdarna (4/4)
talen (2/2)
ställe (9/9)
sekajäte (1/1)
heltidsarbete (2/2)
stiftar (1/1)
husfinska (2/2)
ansiotulo (1/1)
arbetspensionsutdragfinska (1/1)
rörlighet (3/3)
serviceboende (12/12)
App (1/1)
studentbostad (2/2)
Yrittäjän (1/1)
Olkkari (1/1)
undervisning (43/43)
valet (3/3)
utesluta (1/1)
avled (1/1)
blind (1/1)
tillverkning (1/1)
inkassokostnader (1/1)
granskningar (1/1)
utveckla (12/12)
inhämta (4/4)
områdeskoordinatorerna (1/1)
seniorineuvonta (2/2)
brådskande (27/27)
undertecknade (1/1)
fastän (5/5)
handikappet (1/1)
Loktorget (2/2)
kost (2/2)
plats (26/26)
planering (2/2)
ungdomar (27/27)
kredituppgifterna (1/1)
separata (4/4)
torgsidan (1/1)
lähikoulu (1/1)
stipendium (4/4)
strategier (1/1)
ansökningstider (2/2)
tandhälsan (1/1)
fyra (26/26)
läggas (1/1)
försök (1/1)
naturen (11/11)
landets (6/6)
kontakttolkcentral (1/1)
republiken (1/1)
administrerar (1/1)
bolagsmän (1/1)
rekrytering (1/1)
ekonomisk (1/1)
råkar (7/7)
Lahtis (1/1)
dagpenningenfinska (1/1)
underhållsbidraget (4/4)
läsåret (2/2)
bokföring (1/1)
nationalitet (9/9)
bara (13/13)
pedagogiskt (1/1)
upphovsmannens (1/1)
brett (1/1)
personaltjänsteföretag (1/1)
påverkafinska (3/3)
bestämma (10/10)
modersmålsundervisning (1/1)
likvärdiga (2/2)
köper (13/13)
förutsätter (5/5)
könssjukdomarfinska (1/1)
långa (6/6)
tillnyktrings- (1/1)
vokabulär- (1/1)
stadgar (1/1)
ons (3/3)
testamente (5/5)
verkstäder (1/1)
självständighetsdag (1/1)
kartläggning (17/17)
Välkommen (1/1)
grannskapet (1/1)
variera (4/4)
miljötjänster (1/1)
Danske (1/1)
skolanfinska (2/2)
hälsovård (3/3)
nivåer (7/7)
anställdas (5/5)
bott (22/22)
Rösa (1/1)
planera (2/2)
utmärkta (1/1)
vittnen (4/4)
vägra (7/7)
motionsrutter (1/1)
grupplivförsäkring (1/1)
minimilöner (4/4)
finansieras (1/1)
huvudsakligen (2/2)
sistone (1/1)
Sveaborgsfärjorna (2/2)
läroinrättning (2/2)
pdf (25/26) PDF (1)
verksamhetfinska (3/3)
EU- (6/6)
samkönade (2/2)
barnlöshetspolikliniken (1/1)
förlängs (3/3)
förhandsmeddelande (1/1)
riksdag (1/1)
omkring (1/1)
bristfälliga (1/1)
familjerådgivning (5/5)
hoppat (1/1)
missbruksfrågor (1/1)
löpning (1/1)
originalexemplaren (5/5)
grannkommuner (1/1)
från (235/235)
statens (9/9)
utvisningfinska (1/1)
skriftliga (5/5)
Psykologiförbund (1/1)
valmentava (1/1)
toimintaohjelma (1/1)
tukiasuminen (1/1)
skattekortet (6/6)
friluftsmuseum (1/1)
upplysningar (2/2)
juridiska (6/6)
företagarguider (1/1)
skillnad (1/1)
kontakttolkar (1/1)
föds (18/18)
sluta (6/6)
symboler (1/1)
grupperna (1/1)
invånare (45/45)
midsommartraditionerna (1/1)
värms (1/1)
bostadsbidraget (3/3)
där (110/110)
understöd (10/10)
förtroendemannen (4/4)
värdegrunden (1/1)
upphovsrättsavgifter (1/1)
mest (3/3)
mentalvårdsenheten (1/1)
sjunga (2/2)
filmfestivaler (2/2)
Grankulla (40/40)
inbringar (2/2)
krigsskadestånd (1/1)
lokalförvaltning (3/3)
dina (112/113) Dina (1)
Nokia (1/1)
rättegången (2/2)
slussa (1/1)
regent (1/1)
tvingas (5/5)
främja (9/9)
intersexuella (1/1)
make (27/27)
beslutar (13/13)
somrarna (1/1)
bokföringsskyldighet (1/1)
rätten (11/11)
vakuus (1/1)
kvotflyktingens (1/1)
ortodox (4/4)
naturhistoriska (1/1)
Kitfinska (1/1)
föräldrarfinska (1/1)
deltar (6/6)
nationalmuseum (1/1)
norrsken (3/3)
valmansförening (1/1)
Nöteborgsfreden (1/1)
terrängen (1/1)
nämn (1/1)
kreditupplysningsregistret (2/2)
äktenskapet (29/29)
kännas (1/1)
mottagningen (5/5)
privatsektorn (1/1)
händelser (5/5)
bidraget (2/2)
tryggad (3/3)
Jönsasvägen (1/1)
underhyresgäst (3/3)
musikskolorna (1/1)
Steinerskola (2/2)
gymnasie- (1/1)
förföljelse (2/2)
måltiden (1/1)
ett (963/965) Ett (2)
psykiatrisk (2/2)
familjefrågor (4/4)
arbetslöshetstförmån (1/1)
Soites (4/4)
Medelhavet (1/1)
alkoholism (1/1)
finskafinska (2/2)
fungera (2/2)
Centralförbund (1/2) centralförbund (1)
packas (2/2)
tandkliniken (3/3)
studentteaters (1/1)
bifoga (7/7)
sjöstad (1/1)
ekonomibranschen (2/2)
stödmottagarens (1/1)
anmäl (2/2)
socialskyddsförmånerna (1/1)
stadiet (6/6)
pensionspremierna (1/1)
höghusfinska (1/1)
hen (28/28)
arbetarna (2/2)
rekommenderas (2/2)
högskola (7/7)
kontrollerar (1/1)
lagligt (5/5)
treårig (1/1)
Sovjetunionen (8/8)
lärande (4/4)
midsommaren (1/1)
barnförhöjning (1/1)
tidsbeställningfinska (1/1)
upplöses (1/1)
islam (1/1)
persons (3/3)
utövat (2/2)
posttraumatiskt (2/2)
gravplats (1/1)
vanhempainvapaa (1/1)
avfallshanteringfinska (1/1)
nordlig (1/1)
bostadslösas (1/1)
flyktingarna (2/2)
delbeslut (3/3)
kartor (1/1)
månatligen (2/2)
företagstjänsterna (1/1)
förhandsröstningstiden (1/1)
skattefriheten (1/1)
lättläst (1/1)
komma (53/53)
Veroprosentti (1/1)
enspråkiga (2/2)
skattas (1/1)
spalt (1/1)
medborgarefinska (11/11)
kosthålls- (2/2)
examensnivåerna (1/1)
tvingades (1/1)
himmelsfärdsdag (1/1)
lektioner (2/2)
handelsläroanstalten (1/1)
hemvårdens (5/5)
musikinstitutet (1/1)
engelska (783/783)
viktigare (1/1)
studentexamenfinska (1/1)
städerna (7/7)
kom (18/18)
självständighetens (1/1)
arbetsplatserfinska (1/1)
språkinlärning (1/1)
tillräckligt (25/25)
kulturproducenter (1/1)
telefoner (1/1)
ifyllda (3/3)
barnatillsyningsmännen (1/1)
socialarbete (6/6)
möjlighet (23/23)
skuld (1/1)
anmäla (40/40)
tandklinikerna (1/1)
åriga (10/10)
värd (1/1)
ansökningspraxis (1/1)
Danmark (1/1)
balansera (1/1)
varorna (1/1)
legaliseras (4/4)
samboende (1/1)
tidsgränser (1/1)
neuvontapalvelu (1/1)
ovannämnda (1/1)
uppehållstillståndskortet (1/1)
brev (5/5)
anledningarna (1/1)
lönenivån (1/1)
mentorprogram (1/1)
kommunalvalet (2/2)
hyresavtalet (16/16)
ser (8/8)
wc (1/1)
babyresa (1/1)
svartsjuka (1/1)
appar (2/2)
ärendehantering (2/2)
lärare (4/4)
ordnas (81/81)
FIRST (1/1)
avtalats (2/2)
praktiska (7/7)
rederiverksamheten (1/1)
upprättar (3/3)
hörselskada (3/3)
bosniska (2/2)
matburkar (1/1)
service (2/3) Service (1)
bostadsaktier (1/1)
företagarnas (6/6)
erforderliga (1/1)
förstår (1/1)
inbyggd (1/1)
avläggas (5/5)
FPA:s (55/57) Fpa:s (2)
allmänläkare (3/3)
gjorde (1/1)
samtycker (2/2)
saker (27/27)
sammanhang (2/2)
försäljning (1/1)
anslutningsledning (1/1)
bioavfall (2/2)
arbetsavtalet (15/15)
myndighets (1/1)
arbetsförmögen (1/1)
centraler (1/1)
vill (149/149)
jouren (6/6)
socialtjänster (4/4)
priserna (5/5)
ungdomstjänster (6/6)
ställa (6/6)
fiskeområden (1/1)
S2 (4/4)
en (1442/1442)
maj (1/1)
motionera (1/1)
framförd (1/1)
foto (1/1)
työntekijä (1/1)
yöpäivystys (2/2)
sjukskötare (6/6)
densamma (1/1)
Adolf (1/1)
positiva (1/1)
väderförhållanden (1/1)
investerat (1/1)
trakasserier (2/2)
småbarn (1/1)
människohandelfinska (1/1)
HOAS (8/8)
studietakt (1/1)
faktureringstjänst (1/1)
chef (8/8)
frivillig (5/5)
familj (22/22)
föbund (1/1)
verovelvollisen (1/1)
studentrabatter (1/1)
ry:s (2/2)
inkomsterna (6/6)
motionsmöjligheter (2/2)
knapp (1/1)
gardet (1/1)
praktiskt (1/1)
kvar (10/10)
tillhandahålls (9/9)
jobbsökande (2/2)
föräldradagpenningar (3/3)
innefattar (1/1)
kallelsen (1/1)
fortsättningen (1/1)
släktingar (9/9)
tvillingar (1/1)
diplomi (1/1)
bolagsman (2/2)
tillfälliga (3/3)
umgängesrätt (6/6)
luggas (1/1)
ingång (3/3)
lönesättning (1/1)
rutterna (1/1)
musiikkiopisto (1/1)
vårdkostnaderna (1/1)
giftermål (1/1)
pendlar (1/1)
upphängningsbygel (1/1)
integrationsprocessen (1/1)
i (2699/2701) I (2)
tandkliniker (4/4)
invandrarförening (1/1)
modersmål (35/35)
motionshobbyer (1/1)
uppfyllas (1/1)
företagarkurser (1/1)
pensionsförsäkring (3/3)
några (24/24)
tretton (1/1)
notarius (1/1)
skattekort (20/20)
indriver (1/1)
päiväkoti (2/2)
Tölö (2/2)
yngre (5/5)
pitkä (1/1)
jobbsökningen (11/11)
idrottscentret (1/1)
årskurs (5/5)
Uleåborgs (1/1)
kvällarna (1/1)
rutten (1/1)
slutliga (3/3)
siffror (1/1)
utbilda (5/5)
Duo (1/1)
öppningsoperation (3/3)
förstå (2/2)
medborgarinstitutet (1/1)
fattats (4/4)
gentemot (2/2)
automat (1/1)
ytmaterial (1/1)
släktning (1/1)
järnvägsstation (1/1)
bokbussarna (1/1)
EHIC (1/1)
smärtan (1/1)
inredning (1/1)
ge (23/23)
näringsbyråeran (1/1)
klä (4/4)
fackman (1/1)
museidagen (1/1)
Brottsofferjouren (4/5) brottsofferjouren (1)
samfällighets (3/3)
sjöss (3/3)
SOA (1/1)
tillväga (1/1)
barns (19/23) Barns (4)
keskus (1/1)
Gloet (2/2)
mera (5/5)
permanent (17/17)
aktörer (1/1)
ligger (22/22)
idrottsföreningar (1/1)
visumets (1/1)
brottsoffer (1/1)
almanacksbyrå (2/2)
bredvid (1/1)
Celia (1/1)
Rosatom (1/1)
webbutik (1/1)
resepti (1/1)
rättigheterfinska (1/1)
lönsamheten (1/1)
ägarbostäderfinska (2/2)
högskolors (1/1)
religionsfrihet (2/2)
mödrarådgivningstjänsterna (1/1)
hyresgäst (1/1)
omskärelsen (2/2)
gav (2/2)
praktiknära (2/2)
reaali (1/1)
språkversionerna (2/2)
bevittnat (1/1)
försäkringspremierna (4/4)
avlyssnas (1/1)
stämma (3/3)
religiös (5/5)
juridiskt (2/2)
skidåkningfinska (1/1)
avfallsåtervinningfinska (1/1)
kontaktuppgifterna (15/15)
oklarheter (3/3)
onsdagar (4/4)
flyga (1/1)
paluun (1/1)
brottmålet (1/1)
båtliv (1/1)
svensk (1/1)
Pensionsskyddscentralen (6/6)
följa (19/19)
handikapptolkar (1/1)
avgifter (5/5)
ägarskapet (1/1)
godtagbar (3/3)
kursutbudet (1/1)
förvaltas (1/1)
Väestöliittos (2/2)
motionslokaler (1/1)
vigslar (2/2)
remixa (1/1)
vardera (2/2)
kulturell (1/1)
Korso (3/3)
anställningsoptioner (1/1)
frågor (51/51)
enas (2/2)
vikt (1/1)
uppsägningstid (2/2)
toimeentulotuki (1/1)
radhus (3/3)
grundinformation (1/1)
besiktigas (1/1)
parförhållande (24/24)
hjälp (183/183)
ogift (3/3)
Hanhikivi (1/1)
letade (1/1)
utgångstid (1/1)
frånluftsventilerna (1/1)
par (17/17)
trästadshelheter (1/1)
skriftligt (27/27)
utvecklingsstörda (3/3)
situationer (32/32)
plast (1/1)
lönen (16/16)
skolhälsovårdenfinska (1/1)
beställa (14/14)
ingått (6/6)
uppsägning (4/4)
undertecknar (4/4)
umgängesarrangemanget (1/1)
skedda (1/1)
affärsverksamhetsplanen (5/5)
vilka (37/37)
Ryssland (9/9)
antingen (35/35)
paus (1/1)
äitiyspakkaus (1/1)
avger (1/1)
avbryta (2/2)
underhållsbidrag (8/8)
profil (2/2)
läkemedelskostnaderna (1/1)
inkomst (12/12)
handikappad (4/4)
administrativa (2/2)
Barnskydd (1/1)
sekretessplikt (2/2)
förväntar (5/5)
invaliditet (1/1)
upplagan (1/1)
talas (8/8)
läkartid (4/4)
resekostnader (1/1)
slussar (1/1)
leverans- (1/1)
farliga (2/2)
inga (9/9)
högtidlig (1/1)
skolarbete (1/1)
väestötietojärjestelmä (1/1)
mentalvårdstjänster (2/2)
likvärdigt (4/4)
främjar (5/5)
ut (113/113)
visar (2/2)
försäkringen (4/4)
fiskebyn (1/1)
portfölj (1/1)
form (11/11)
Israel (1/1)
slottfinska (1/1)
utbildningsprogrammen (2/2)
stödnät (1/1)
matkakortti (2/2)
Unionin (1/1)
sysslorna (3/3)
fysiska (4/4)
upptagna (1/1)
hyrestiden (3/3)
högskoleutbildning (5/5)
äldre- (1/1)
våldssituationer (1/1)
markområden (1/1)
långt (4/4)
metspö (3/3)
sambor (5/5)
kuntoutuspäätös (1/1)
Lapin (1/1)
verkställer (1/1)
Tallinn (2/2)
känslofyllda (1/1)
bolag (6/6)
erövrade (2/2)
hjälpa (26/26)
matkulturenengelska (1/1)
tvätten (1/1)
socialhandledarna (1/1)
lähdevero (1/1)
klinikka (3/3)
elapparater (1/1)
papper (5/5)
backe (1/1)
valt (1/1)
vårda (1/1)
årskurserna (12/12)
årstider (2/2)
käyttövastike (1/1)
professionella (1/1)
hyresavtal (16/18) Hyresavtal (2)
rummet (1/1)
metall (1/1)
studerandeengelska (1/1)
bil (12/12)
perintövero (1/1)
kompetens (3/3)
nog (1/1)
byggas (1/1)
Rinteenkulma (1/1)
diskuteras (1/1)
hyrorna (1/1)
bastulaven (1/1)
företag (101/101)
vuxenstuderande (4/4)
Förenta (1/1)
tjänst (11/11)
teckenspråketfinska (1/1)
repertoar (1/1)
forskningen (1/1)
tryggaste (2/2)
aikuisopisto (6/7) Aikuisopisto (1)
inleder (6/6)
ungdomsarbete (3/3)
t.ex. (18/18)
antagning (1/1)
remiss (12/12)
värde (1/1)
regioner (1/1)
telefonnummer (8/8)
informellt (1/1)
preventivmedels- (1/1)
särskilda (5/5)
grenarna (1/1)
tvåspråkighet (1/1)
framställningen (2/2)
matsäck (1/1)
jobbar (1/1)
sökningen (1/1)
Takuusäätiös (1/1)
överhuvudtaget (1/1)
kommunalt (3/3)
plastprodukter (2/2)
anordnas (5/5)
hjälpt (1/1)
arbetslöshetsförmån (7/7)
integrationen (4/4)
bostadsrättsbostaden (1/1)
spelar (1/1)
www.gramex.fi (1/1)
verklig (2/2)
åldringspension (1/1)
förutsätta (1/1)
kaksoistutkinto (1/1)
människovärde (1/1)
skarvsladd (1/1)
skatterelaterade (1/1)
livsåskådning (1/1)
upprättade (1/1)
Versofinska (1/1)
universitets- (1/1)
kemiska (1/1)
apoteket (8/8)
dator (5/5)
förvärvar (1/1)
bekymrar (1/1)
utsända (1/1)
reseplaneraren (3/5) Reseplaneraren (2)
tingsrätten (9/9)
dagvårdsplatsen (1/1)
undersökningarna (5/5)
huvudbiblioteket (1/1)
fackets (1/1)
mamman (1/1)
upprätthåll (1/1)
makarnas (6/6)
fullgjort (1/1)
kvinna (3/3)
intervjuer (1/1)
utrikesministeriet (2/2)
medicinska (2/2)
tillämpas (6/6)
undantag (4/5) Undantag (1)
företagaren (5/5)
socialnämnden (1/1)
Flyktingrådgivningens (1/1)
motionsslingor (3/3)
pensionsåldern (1/1)
ansvarsområden (1/1)
allmänna (18/18)
osäker (2/2)
försenad (2/2)
avvisa (2/2)
tysta (4/4)
yrkesläroanstalterfinska (1/1)
kropps (1/1)
mamma (1/1)
telegram (1/1)
ansökan (145/147) Ansökan (2)
tips (3/3)
invandrarenheten (2/2)
politiskt (1/1)
smarta (1/1)
jämställdhet (12/14) Jämställdhet (2)
beroende (10/10)
ställer (2/2)
förutom (2/2)
behörig (1/1)
nedtecknas (2/2)
pensioner (2/2)
skoltiden (1/1)
rabatt (5/5)
sommaren (10/10)
styrgrupp (1/1)
bifaller (1/1)
överstiga (2/2)
notaries (1/1)
mellan (40/40)
brandvarnare (6/6)
ordnades (1/1)
studietiden (1/1)
Flyktingrådgivningen (3/3)
befogad (1/1)
kvinnorfinska (1/1)
förvaltning (1/1)
arbetskraftsutbildning (18/19) Arbetskraftsutbildning (1)
mellannivån (1/1)
sjöfartsbranschen (1/1)
förberedelserna (2/2)
vårdledighet (4/4)
biografens (1/1)
han (44/44)
datorn (1/1)
öster (2/2)
hälsovårdarens (3/3)
mottagningar (2/2)
handikappråd (1/1)
yrkeskunnighet (7/7)
framföra (2/2)
undrar (1/1)
förskoleundervisning (14/15) Förskoleundervisning (1)
yrkesprov (1/1)
kommunallagen (1/1)
inletts (1/1)
Havukoski (1/1)
ny (12/12)
undervisningstimmar (1/1)
basis (11/11)
återkallas (6/6)
föreningar (13/14) Föreningar (1)
specialdiakoner (1/1)
mannen (5/5)
registerstryrelsen (1/1)
företagsekonomiska (1/1)
Lastensuojelulaki (1/1)
webbläsare (1/1)
rättvisa (1/1)
medicinerna (1/1)
konstaterar (1/1)
beskattningsbeslutet (4/4)
värden (1/1)
handläggningsavgiften (1/1)
ensam (15/15)
campingområdenfinska (1/1)
vakinaista (2/2)
arbetslösheten (4/4)
lunchpaus (1/1)
energiavfall (2/2)
verifierats (1/1)
hälsomyndighet (1/1)
förmånligaste (1/1)
PB (1/1)
tjänstemän (1/1)
Liitto (4/4)
fullföljer (1/1)
varainsiirtovero (1/1)
stängd (1/1)
beskriva (1/1)
toisena (1/1)
två (97/97)
genomgått (1/1)
koncernen (1/1)
samboförhållande (14/16) Samboförhållande (2)
räntorna (1/1)
bekosta (3/3)
stödtjänsterfinska (1/1)
äldsta (2/2)
företer (1/1)
skilsmässafinska (2/2)
samkommunens (1/1)
utföras (3/3)
stödperson (4/4)
grundandet (1/1)
videon (1/1)
startar (5/5)
forskarefinska (1/1)
bilplats (1/1)
revisionsbyråer (1/1)
Internetberoende (1/1)
ansökningen (7/7)
hjälper (63/63)
etnisk (2/2)
Yle (1/1)
metalli (1/1)
republik (2/2)
matlagning (3/3)
bättre (5/5)
rehabiliteringen (5/5)
genomgå (2/2)
kontorenfinska (1/1)
Schengenland (1/1)
informationstjänst (1/1)
Fennovoimas (1/1)
lär (16/16)
vårdenheter (1/1)
å (3/3)
samfunden (1/1)
fyllt (29/29)
prepaid (2/2)
CVfinska (2/2)
betalningspåminnelse (1/1)
Studieinfo.fi (9/9)
direktör (1/1)
inleda (3/3)
köpa (32/33) Köpa (1)
taxin (1/1)
kollektivtrafiken (4/4)
priset (2/2)
tolkförbunds (1/1)
magistrat (4/4)
tillgångar (4/4)
sammanlagda (2/2)
förhöjd (1/1)
stadenfinska (3/3)
postadressen (1/1)
namnskylt (1/1)
flaggdagarna (1/1)
droganvändning (1/1)
arbetslagstiftningenfinska (1/1)
köra (6/6)
försäkringarna (1/1)
kommunstyrelsen (1/1)
kymppiluokka (2/2)
uppstartsföretagarefinska (1/1)
danska (2/2)
webbplats (174/174)
työehtosopimukset (1/1)
hjälpsystemet (1/1)
betyder (24/24)
språkfinska (2/2)
arvsskattfinska (1/1)
inresa (1/1)
likabehandling (12/12)
uppfostrande (1/1)
gäster (1/1)
klassen (4/4)
december (6/6)
HIVfinska (1/1)
finansrådgivningen (1/1)
polisanmälan (1/1)
könen (2/2)
servicerådgivningen (1/1)
sätt (44/44)
karttjänstfinska (1/1)
välfungerande (1/1)
läroplikten (2/2)
använder (17/17)
työtulo (1/1)
paperi (1/1)
handikapptjänsternafinska (1/1)
muntligt (2/2)
museum (3/3)
Esbo (100/100)
ängarna (1/1)
ungdomsledare (1/1)
Esbotillägget (1/1)
työvoimakoulutus (1/1)
märker (1/1)
avgångsbetyget (1/1)
vardagssysslor (2/2)
specialundervisningen (1/1)
bildar (1/1)
rätt (226/226)
jakttillstånd (1/1)
länkarna (2/2)
examen (68/68)
ungafinska (8/8)
video (2/2)
upplever (7/7)
gåva (1/1)
förseningsavgift (1/1)
försenade (2/2)
bokad (1/1)
besitter (1/1)
förekommer (2/2)
familjemedlemmen (1/1)
studieprogrammet (1/1)
skolpsykologerna (1/1)
livsmedel (2/2)
antagits (2/2)
efternamnfinska (1/1)
lyssna (2/2)
ställt (2/2)
makar (2/2)
områdena (1/1)
skaffar (6/6)
sopkärlen (1/1)
betjänad (1/1)
ovanliga (1/1)
uppväxt (4/4)
socialarbetarefinska (1/1)
helhetsbetonade (1/1)
handledning (21/21)
borgerlig (2/2)
frivilligarbete (5/6) Frivilligarbete (1)
kurator (1/1)
beviljar (4/4)
hälsovårdsbranschen (1/1)
karttjänsten (2/2)
Veikko (1/1)
handelsregisterutdraget (1/1)
principerna (1/1)
renoveringskostnaden (1/1)
fryser (1/1)
flexibla (1/1)
trafikerar (1/1)
språket (50/50)
plastleksaker (1/1)
stödcentretfinska (1/1)
självrisk (1/1)
orterna (1/1)
de (328/335) De (7)
boendemöjligheter (1/1)
hämtas (1/1)
grundats (2/2)
ångest (1/1)
Rovaniemiområdet (1/1)
bostadsaktiebolagets (2/2)
pompa (1/1)
noggrann (2/2)
senioruniversitetet (2/2)
begått (4/4)
förhållande (1/1)
ITE (1/1)
ansökt (4/4)
missnöjd (1/1)
obligatoriska (4/4)
lön (46/46)
aurora (1/1)
honom (3/3)
Tavataan (1/1)
färdighetsnivåerna (1/1)
verksamhetsprogram (1/1)
organisationerna (1/1)
rubriken (8/8)
förpliktelser (1/1)
resurser (2/2)
specialtillstånd (1/1)
matställen (1/1)
Liikenteen (1/1)
invånarparker (1/2) Invånarparker (1)
jourtid (1/1)
bemärkelsedagar (1/1)
statligt (1/1)
ålderfinska (1/1)
legalisera (1/1)
dagsgymnasierna (1/1)
kierratys.info (2/2)
tillståndsansökningarfinska (1/1)
serbiska (1/1)
vardagar (17/17)
elpriserfinska (1/1)
isolering (1/1)
stämman (1/1)
omfattar (24/24)
utbytesstudenter (1/1)
ersättningarfinska (1/1)
bostadsrådgivning (1/1)
kliniken (7/8) Kliniken (1)
skattskyldiga (1/1)
rusmedels- (1/1)
munsjukdomar (1/1)
finsk (51/51)
särbehandlas (2/2)
rörelsehindradefinska (1/1)
klinikerna (1/1)
karens (1/1)
fortsatta (9/9)
invandrarungdomar (1/1)
pensionen (2/2)
nytt (26/26)
menar (1/1)
registreringsblanketten (1/1)
idrottshallar (2/2)
rådgivningsbyrå (2/2)
högsta (8/8)
Card (1/1)
bidrag (11/11)
och (2619/2619)
kyrkor (1/1)
bilen (6/6)
utgången (4/4)
kristelefon (3/3)
asylsökandefinska (2/2)
daghemmet (7/7)
socialväsendet (1/1)
tobaksprodukter (1/1)
släktband (1/1)
stadsmuseum (1/1)
föräldrapenningperiodens (1/1)
ställningen (1/1)
Handikappforums (1/1)
sjukhus (31/31)
känner (12/12)
vila (1/1)
mottagningscentral (4/4)
uppfylls (4/4)
socialtjänst (1/1)
folkhögskolanfinska (1/1)
snöskottande (1/1)
Villenpirtti (1/1)
USA (4/4)
större (13/13)
arbetsmarknadsstöd (4/4)
invandrareleverna (1/1)
linkkiBybiblioteken (1/1)
sociala (74/74)
byggs (1/1)
icke (5/6) Icke (1)
konditionen (2/2)
tog (3/3)
studiefärdigheter (1/1)
startsida (1/1)
initiativ (1/1)
färdtjänst (7/7)
judarna (1/1)
Jorv (10/10)
tillgångarna (1/1)
detsamma (1/1)
varmt (2/2)
betalningsplan (2/2)
barndom (1/1)
Opintopolku.fi (3/3)
Genève- (2/2)
helgjour (1/1)
kistor (1/1)
alkohol- (3/3)
motorfordon (3/3)
avsnitten (1/1)
åsikter (3/3)
riskfaktorer (1/1)
utbildningenfinska (1/1)
användaren (2/2)
företagsläkare (1/1)
missbrukarproblem (2/2)
standardblanketter (1/1)
semestern (2/2)
FPA.Som (1/1)
församlingars (1/1)
blommor (2/2)
olycksfall (5/5)
finska (348/355) Finska (7)
rådgivningens (1/1)
kraftig (1/1)
arv (2/2)
granskas (1/1)
högst (37/37)
vänskap (1/1)
höghus (10/10)
Perheiden (2/2)
fordonsföreskrifter (1/1)
hotad (1/1)
rokotus (1/1)
progressivt (1/1)
medlemmars (2/2)
enkelt (2/2)
finansiera (1/1)
bekräftade (1/1)
sosiaalineuvonta (1/1)
folkhögskolor (3/3)
handläggarna (1/1)
lönesystemet (1/1)
utbildningsprogrammet (1/1)
databas (1/1)
cykla (4/4)
serviceställe (5/5)
närståendevårdfinska (6/6)
stad (47/47)
Röda (10/15) röda (5)
består (8/8)
henne (4/4)
byråns (13/13)
hyr (8/8)
riskabelt (1/1)
avausleikkaus (2/2)
vapaarahoitteinen (1/1)
enbart (3/3)
sommarlov (1/1)
tolktjänsterna (4/4)
teknik (2/2)
stridig (1/1)
befolkningsdataregistret (1/1)
rådgivare (1/1)
flerårigt (1/1)
intervjuerna (1/1)
ettdera (1/1)
skett (1/1)
biblioteketfinska (2/2)
besvärsanvisning (1/1)
orolig (2/2)
träna (1/1)
cycling (1/1)
täckjacka (1/1)
villasamhället (1/1)
villkor (18/18)
hälsostationerna (10/10)
Asuntosäätiös (1/1)
skola (18/18)
byggnader (2/2)
barnets (93/94) Barnets (1)
era (2/2)
patientförening (1/1)
skidspår (2/2)
svarar (6/6)
rehabiliteringfinska (5/5)
isännöitsijä (1/1)
uppgöra (1/1)
avsedda (27/27)
adressen (10/10)
MTV3 (1/1)
aktiebolag (4/4)
påskdagen (1/1)
kvotflyktingarna (1/1)
specialist (6/6)
minderårig (2/2)
ansöker (72/72)
anses (10/10)
festivalerfinska (1/1)
borgarna (1/1)
medelstora (1/1)
assistent (1/1)
könsstympning (2/2)
dari (2/2)
Perho (1/1)
emigranter (2/2)
kundrådgivningen (1/1)
rasismi (1/1)
idrottsanläggningarna (1/1)
osaomistusasunto (2/2)
peruskoulutukseen (1/1)
inkorporerade (1/1)
adresserna (1/1)
tillåtelse (1/1)
Kors (9/11) kors (2)
aktuella (6/6)
angett (1/1)
bosättningsort (1/1)
tel (2/2)
bevisar (2/2)
dubbelrum (1/1)
offentlig (8/8)
ljusa (1/1)
kortvarigt (1/1)
papparollen (1/1)
kotoutumissuunnitelma (1/1)
teatrarnas (2/2)
naturkunskap (1/1)
återgå (3/3)
rullator (1/1)
men (71/71)
projektet (1/1)
sista (6/6)
konstämnen (3/3)
traditionell (2/2)
föreningarna (1/1)
flyktingkvoten (1/1)
syn (2/2)
äktenskapsförord (4/5) Äktenskapsförord (1)
skriftligen (2/2)
individer (1/1)
hem (34/34)
asiointipiste (1/1)
hemma (39/39)
nomineras (2/2)
delegation (1/1)
elektrisk (2/2)
näromgivning (2/2)
advokater (1/1)
familjevåldfinska (2/2)
omedelbart (3/3)
osasairauspäiväraha (1/1)
invandrarkunder (1/1)
Nettineuvola (1/1)
avancemang (2/2)
tand- (1/1)
lägger (2/2)
period (5/5)
republikens (1/1)
egentliga (4/4)
tvingande (2/2)
partiella (3/3)
växte (1/1)
ungdomsgård (2/2)
Finlandengelska (6/6)
grad (1/1)
lönar (17/17)
synnerligen (1/1)
penningunderstöd (2/2)
beredning (2/2)
fullsatta (1/1)
Vantaalla.info (1/1)
skolan (43/43)
språkstudier (1/1)
upprepade (1/1)
koncentrerad (1/1)
gymnasiebaserad (2/2)
fortsättare (1/1)
uppföljning (1/1)
servicehandledaren (1/1)
brandsläckare (1/1)
kränker (1/1)
språkkurserna (1/1)
röstningsställe (1/1)
genom (47/47)
bedriver (5/5)
utsidan (1/1)
kontinuerligt (8/8)
psykologen (2/2)
spelproblem (4/4)
jobbsökningfinska (1/1)
reparationsarbeten (1/1)
vidimeras (1/1)
ske (2/2)
helheter (1/1)
berätta (5/5)
Karlebystödet (1/1)
rötter (1/1)
natur (1/1)
stater (2/2)
tillräckliga (25/25)
gett (2/2)
kontoutdrag (1/1)
förslossningsdatumet (1/1)
personliga (3/3)
underhållet (1/1)
Företagsfinland (1/1)
platsen (1/1)
utbudet (3/3)
underhållsbehov (3/3)
enhetlig (1/1)
otrogenhet (1/1)
betald (1/1)
bostadsform (1/1)
kylskåpet (2/2)
verksamheter (1/1)
forna (1/1)
Björkby (2/2)
misstänks (2/2)
studentkort (1/1)
nedan (1/1)
-motion (1/1)
mödrarådgivning (1/1)
EK (2/3) Ek (1)
motionsalternativfinska (1/1)
valomgången (3/3)
räkna (2/2)
mobbning (1/1)
hemstad (2/2)
terminsavgift (1/1)
skada (8/8)
lutherska (19/19)
växel (1/1)
samlaget (1/1)
itsenäisen (1/1)
situationen (14/14)
museer (10/10)
rådgivnings- (2/2)
trossamfund (5/5)
institutfinska (1/1)
Vanda (115/115)
graviditeten (16/16)
ljudet (1/1)
arvonlisävero (1/1)
fötts (3/3)
bemött (1/1)
näringfinska (1/1)
moderns (7/7)
bindande (6/6)
genomförandet (1/1)
avslutar (1/1)
bransch (9/9)
NewCo (5/5)
pääomatulo (1/1)
Schengen (1/1)
rester (1/1)
möjlig (2/2)
födelsedatumet (1/1)
akutmottagningen (1/1)
socialbyrån (15/15)
sjukvårdsdistrikt (3/3)
drog- (1/1)
bröllopsdagen (1/1)
målsättningar (1/1)
buddhism (1/1)
löneinkomster (2/2)
samarbetet (2/2)
föder (4/4)
helst (23/23)
julens (1/1)
parkera (1/1)
samkommunen (3/3)
bioprogram (1/1)
tidsbokningstjänst (1/1)
förberedande (39/41) Förberedande (2)
aktiviteter (10/10)
lettiska (1/1)
Centralförbundet (1/1)
skadan (2/2)
upprätthåller (4/4)
barnens (7/7)
äitiysraha (2/2)
Tukiliittos (1/1)
självständiga (3/3)
arbetspensionsanstalt (1/1)
Grankullafinska (1/1)
förskott (1/1)
Startpunkter (1/1)
Kela (11/11)
Ohjaamo (1/1)
medeltemperaturen (1/1)
bekräftats (2/2)
samarbetar (1/1)
jourmottagning (1/1)
integrationsrelaterade (4/4)
babyskydd (1/1)
kön (22/22)
vittna (1/1)
området (18/18)
samband (10/10)
tolkförbund (2/2)
saknas (2/2)
sitt (53/53)
agera (1/1)
borde (2/2)
festföremålet (1/1)
garantier (1/1)
FIRMAXI (1/1)
åsikt (8/8)
diskriminera (3/3)
prata (12/12)
utvisning (1/1)
Strandväg (1/1)
dagvård (10/11) Dagvård (1)
Befolkningsregistercentralen (1/1)
sidorna (9/9)
hälsomotionsgrupper (1/1)
familjeförmåner (2/2)
obegränsat (1/1)
oartigt (3/3)
flerfaldiga (1/1)
ansökningens (1/1)
gymnasieutbildningen (1/1)
centralen (2/2)
telefonrådgivning (3/3)
anställningsintervju (1/1)
läcker (1/1)
storindustrin (1/1)
Migrationsverket (28/31) migrationsverket (3)
passa (1/1)
hantverk (3/3)
utkomststöd (18/18)
pappersblankett (5/5)
insjuknade (1/1)
uppskatta (4/4)
linkkiFörbundet (1/1)
diskmaskinen (2/2)
tidigare (21/21)
religionstillhörigheten (1/1)
jämställdheten (1/1)
studieresultat (1/1)
stadinasunnot.fi (1/1)
mån.-tors. (1/1)
fanns (3/3)
tävlingen (4/4)
införd (1/1)
mikrovågsugnen (1/1)
nära (13/13)
ljudböcker (2/2)
skrivas (3/3)
avfall (10/10)
anslutet (2/2)
februari (5/5)
papperspåse (1/1)
trappan (1/1)
beräknade (6/6)
familjemedlemmarna (2/2)
pyssel (1/1)
avgiftsbelagda (9/9)
allvarliga (1/1)
familjeförhållanden (4/4)
förändringsarbeten (2/2)
finskt (30/34) Finskt (4)
straffbart (2/2)
lämnas (13/13)
mödravården (2/2)
yliopisto (4/4)
EU (117/117)
ordningsregler (2/2)
produkter (5/5)
anhörigfinska (1/1)
intjänade (3/3)
kauniainen.fi (1/1)
kulturevenemang (1/1)
stadsbiblioteken (1/1)
rättigheterna (2/2)
kvinnan (5/5)
ganska (1/1)
Omena (4/4)
minoriteter (3/3)
bostadsort (2/2)
vårdledigheten (2/2)
borealis (1/1)
högskolestudier (8/8)
ledare (1/1)
integrationfinska (1/1)
uttalas (1/1)
föräldrar (37/37)
integrera (2/2)
diakoniarbetaren (1/1)
kansliet (1/1)
osakligt (3/3)
Kanada (1/1)
stödåtgärderfinska (1/1)
dokumentmallar (1/1)
allmänt (6/6)
sökandens (2/2)
önskar (5/5)
härsken (1/1)
DVD (1/1)
skicka (27/27)
maken (10/10)
nattetid (1/1)
försvarsmakt (1/1)
rättshjälpsbyrån (4/4)
betalats (3/3)
skåp (1/1)
förmiddagen (1/1)
veta (4/4)
mödrarådgivningen (8/8)
utbildningsstöd (1/1)
kontaktuppgifterfinska (7/7)
sjukdomar (8/8)
acceptansen (1/1)
arbetslöshet (2/2)
on (2/2)
stressyndromfinska (1/1)
högljutt (3/3)
näringsbyråns (9/9)
hushåll (7/7)
cirkus (1/1)
finansieringsandelar (1/1)
kommunernas (4/4)
vårdnadshavares (1/1)
fordrar (1/1)
visumansökan (1/1)
datumet (2/2)
traumatiska (1/1)
skulden (2/2)
leksaker (2/2)
parkeringsautomater (1/1)
vidare (10/10)
universitetsutbildningar (1/1)
konventionerna (2/2)
meddela (18/18)
idkandet (1/1)
Takuusäätiö (3/3)
märkts (1/1)
ca (4/4)
säätiö (1/1)
konfidentiella (2/2)
Opiskelija (4/4)
västliga (1/1)
familjebidrag (1/1)
kopia (4/4)
akutpreventivmedel (1/1)
just (4/4)
närarbetets (1/1)
definieras (4/4)
heltidsarbetande (1/1)
synskada (1/1)
förvärvsinkomster (1/1)
ledande (2/2)
Isyyden (1/1)
någon (71/71)
terapeut (1/1)
företagarens (3/4) Företagarens (1)
jämlika (1/1)
Stenängens (1/1)
busstidtabellerna (1/1)
praxis (1/1)
arbetstagare (32/33) Arbetstagare (1)
lovade (1/1)
ingick (1/1)
VVO (1/2) Vvo (1)
belastad (1/1)
vare (5/5)
skick (7/7)
insamlingsställe (1/1)
regeringenfinska (1/1)
näringsidkare (5/5)
rasism (4/4)
ansökningsblanketter (2/2)
våldsam (3/3)
upprätthålls (5/5)
disponenten (3/3)
våld (57/61) Våld (4)
urval (1/1)
integrationsplaner (1/1)
ansöka (206/206)
varandras (1/1)
hammashoitola (2/2)
resväg (1/1)
sistnämnda (1/1)
tingsrättens (5/5)
riket (1/1)
högskolestuderande (1/1)
anställer (1/1)
aptit (1/1)
uppsikt (3/3)
handredskapsavgiften (1/1)
gymnasiestudierna (2/2)
lånat (1/1)
Myrkytystietokeskus (1/1)
kulturgrupper (1/1)
Kaustarviken (1/1)
uppvisande (1/1)
graviditetsprevention (2/2)
tillfällen (1/1)
endast (44/44)
korrigerande (1/1)
varav (6/6)
nöjaktiga (3/3)
integrering (1/1)
cykelkarta (1/1)
uppskattar (4/4)
cykelvägar (2/2)
staden (32/32)
sairausvakuutus (4/4)
likaså (2/2)
skyldighet (7/7)
engångskaraktär (1/1)
sovittelu (2/2)
uppfyller (5/5)
pappor (1/1)
belönas (1/1)
registrerar (7/7)
tillfrågad (1/1)
arvolaki (1/1)
handleder (8/8)
drogfritt (1/1)
utlandsresa (1/1)
flit (1/1)
muslimska (1/1)
rikt (1/1)
skickar (12/12)
konventioner (1/1)
samtals- (1/1)
sanning (1/1)
hemland (20/20)
servicen (1/1)
fackförbund (14/16) Fackförbund (2)
rådgivningsbyrån (21/21)
medborgarinstituten (1/1)
befinner (5/5)
unga (72/72)
Finlex (2/2)
IT (1/1)
sagotimmar (1/1)
Esbofinska (3/3)
övningsskola (1/1)
Hilma (1/1)
göra (73/73)
Hörselförbundetfinska (1/1)
hos (167/167)
vaccinationer (4/4)
Hollihaan (1/1)
mars (6/6)
Valvira (3/3)
omständigheterna (1/1)
officiell (4/4)
söder (1/1)
man (251/251)
hemresan (2/2)
genomför (1/1)
fortsätter (2/2)
examenfinska (1/1)
gemensam (8/8)
allt (17/17)
utförande (1/1)
glasförpackningar (1/1)
elbolaget (1/1)
betjänar (29/29)
tvåspråkig (1/1)
återresa (2/2)
kielikahvila (1/1)
psykolog (3/3)
Suomi (1/2) suomi (1)
telefontjänster (1/1)
kontinuerlig (1/1)
kaavinta (1/1)
översatt (2/2)
universiteten (3/3)
timmarna (1/1)
medborgarinstitutets (4/4)
yrkesutbildningfinska (4/4)
baserad (2/2)
missbruksproblem (6/7) Missbruksproblem (1)
presidenten (3/3)
röstar (2/2)
tal (1/1)
beskattas (2/2)
inbördeskrig (1/1)
mödrarådgivningar (1/1)
förutsättning (1/1)
förtrogna (1/1)
avvägs (1/1)
kostnadsersättningfinska (1/1)
affärsmodell (1/1)
ställen (3/3)
biblioteken (6/6)
tydliga (1/1)
familjehem (2/2)
arbetsoförmögen (2/2)
bekräftar (5/5)
romerna (1/1)
privatskola (2/2)
representant (2/2)
flyttgodsfinska (1/1)
resedokument (3/3)
bo (55/55)
sälfångst (1/1)
finskundervisning (2/2)
belägna (3/3)
juli (7/7)
flyktingar (14/14)
kronologisk (2/2)
internationalisering (1/1)
pakolainen (1/1)
insamlingskärl (2/2)
bostadsförmedlingar (1/1)
husets (8/8)
läge (1/1)
yrkeskunskaper (2/2)
farförälder (2/2)
ljud (1/1)
föräldrapenningperioden (3/3)
allvarligt (4/4)
fester (3/3)
Seremoniat (1/1)
annat (135/135)
integrations- (2/2)
bildats (2/2)
näringsbyråer (2/2)
kartläggningar (1/1)
gammalt (6/6)
ulosotto (1/1)
förmedlingsarvode (1/1)
dagars (1/1)
polisens (8/9) Polisens (1)
akutvården (1/1)
oljevärme (1/1)
närliggande (2/2)
skolbarn (2/2)
ris (1/1)
kortfattad (1/1)
utbetald (1/1)
ens (3/3)
apotek (4/4)
Nimettömät (1/1)
socialskyddsförmåner (1/1)
flytthjälp (1/1)
boendeservice (2/2)
brinna (3/3)
monteringsarbetsplats (1/1)
kommunikationskanal (1/1)
näst (1/1)
familjeförhållandena (1/1)
öppning (1/1)
beviljats (11/11)
arktiska (3/3)
skärgård (1/1)
studiepoäng (2/2)
studierna (26/26)
dvs. (3/3)
verkar (2/2)
veckoslut (15/15)
barnkapning (1/1)
rehabiliteringscenter (1/1)
stödbostad (3/3)
lika (15/15)
verksamheten (14/14)
barnskyddfinska (1/1)
työpaikat (2/2)
tätorterna (1/1)
därför (5/5)
födelsedagar (1/1)
släktens (1/1)
Tullrådgivningen (1/1)
arbetarskyddsmyndigheterna (3/3)
utbildningarfinska (2/2)
prevention (5/5)
oberoende (5/5)
påfrestande (2/2)
scenkonst (1/1)
församlingens (1/1)
Seure (1/1)
rehabiliteringsbehovet (1/1)
narkotika (1/1)
RIKU (1/1)
förskottsinnehållning (2/2)
runt (29/29)
telefonen (2/2)
vidaredistribuera (1/1)
förtida (3/3)
grunderfinska (1/1)
populär (1/1)
vi (11/15) Vi (4)
väderleksrapporterna (1/1)
magistraternafinska (1/1)
visas (5/5)
alltså (25/25)
tryckta (1/1)
anmärkning (2/2)
hotfullt (1/1)
våldet (1/1)
Finlands (67/67)
driva (5/5)
studentmössor (1/1)
talar (6/6)
depression (2/2)
ympärileikkaus (3/3)
julafton (2/2)
hjälpen (8/8)
tvätta (2/2)
idag (2/2)
serviceplanen (1/1)
handel (1/1)
nättjänsten (2/2)
klasser (5/5)
statsrådet (2/2)
avsett (10/10)
medlemskommuner (1/1)
sparat (1/1)
barnomsorgen (1/1)
rahoitusvastike (1/1)
Määräaikainen (1/1)
ges (42/42)
Kehitysvammaisten (1/1)
MoniNet (4/4)
Wien (2/2)
salu (3/3)
talous- (1/1)
samarbeta (1/1)
sosiaalivirasto (1/1)
läkarutlåtande (2/2)
fastlagsbullar (1/1)
frilansarefinska (1/1)
handikapporganisationer (1/1)
rehabiliteringstjänster (1/1)
köping (1/1)
seglare (1/1)
lyder (1/1)
behov (38/38)
händelsen (1/1)
uskonnonvapaus (1/1)
löneutbetalningen (4/4)
hävs (1/1)
arabisktalande (1/1)
Finnkinos (1/1)
kölapp (1/1)
utreda (5/5)
pojken (2/2)
hälsovårdssamkommun (7/7)
Konsumentförbunds (1/1)
utifrån (10/10)
arbetsplatsintroduktion (1/1)
hobbystudier (2/2)
verben (1/1)
arbetslivetfinska (1/1)
ABC (2/2)
såsom (23/23)
yrittäjien (1/1)
lähityön (1/1)
högskolexamen (1/1)
förlängning (2/2)
ända (3/3)
framsteg (1/1)
dela (5/5)
arbetsgivarna (4/4)
tvätt (1/1)
medier (3/4) Medier (1)
snitt (1/1)
Köpcentret (1/1)
personligt (6/6)
umgänget (4/4)
äitiysneuvola (2/2)
Ludvig (1/1)
arbetslösafinska (3/3)
låneräntan (1/1)
hemlika (1/1)
publicerats (3/3)
Clinic:s (1/1)
förskottsuppbördsregister (1/1)
partiellt (2/2)
friluftsområden (1/1)
utgör (2/2)
fornlämningsområde (1/1)
mandatperioder (1/1)
huvudstad (3/3)
serbokroatiska (1/1)
undervisningsspråket (7/7)
bekräftas (1/1)
delaktighet (1/1)
musikhobby (1/1)
kommunsidor (1/1)
kommunikationsteknik (1/1)
ändamålet (1/1)
studieplats (29/29)
personbeskattning (1/1)
bönder (1/1)
översätta (1/1)
företagsledning (1/1)
bostadslösa (5/5)
kvotflyktingarfinska (1/1)
kommunsida (1/1)
köksskåpen (1/1)
Schengenländer (1/1)
E303 (1/1)
Europaparlamentsvalfinska (1/1)
licentiatexamen (1/1)
perheneuvola (6/6)
dömas (5/5)
Företagarna (1/1)
filmfestival (1/1)
billigaste (1/1)
närvara (1/1)
känns (1/1)
städning (1/1)
ljust (1/1)
YEL (1/1)
skrämma (1/1)
anställningens (3/3)
vintersporterna (1/1)
arbetspraktik (3/3)
titta (5/5)
samtala (2/2)
bevis (4/4)
Suomipassi (1/1)
arbetspensionsanstalter (1/1)
kortvariga (2/2)
slutarbete (2/2)
förlängas (3/3)
tjänsteställen (1/1)
bygger (1/1)
jäte (1/1)
gymnasier (6/6)
annars (5/5)
dagstidning (1/1)
hemsidorfinska (1/1)
bostadsrättsavtal (1/1)
tolktjänster (5/5)
undantagsfall (4/4)
erfarenheter (3/3)
töms (1/1)
seniorer (6/6)
huvudstadsregionens (3/3)
anmälan (25/25)
utgöra (4/4)
huvuddukar (1/1)
är (1322/1322)
teckenspråk (3/3)
expertråd (1/1)
veckor (12/12)
äktenskapsförordet (2/2)
yrkenfinska (1/1)
gränserna (2/2)
återvinningsstation (1/1)
morgonen (7/7)
arbetsmotivation (1/1)
båtlivfinska (1/1)
motsvarar (11/11)
läraren (3/3)
anslöts (2/2)
raskauden (1/1)
Petäjävesi (1/1)
terapeuten (1/1)
fakturor (1/1)
pålitlig (3/3)
användningsdatumet (1/1)
väldigt (4/4)
mellanrum (4/4)
Myyrinkis (1/1)
arbetslivsfärdigheter (2/2)
sjukvårdskortetfinska (2/2)
studenthem (1/1)
stöttar (1/1)
varar (20/20)
levnadskostnader (2/2)
vrida (1/1)
förtrogen (1/1)
överenskommit (1/1)
slutexamen (1/1)
utbildningsplats (2/2)
meddelandet (2/2)
reglerat (4/4)
målet (4/4)
gymnasieelever (1/1)
tohtori (1/1)
påvisa (3/3)
lyfter (1/1)
bevisa (6/6)
Avara (2/2)
advokatförbund (1/2) Advokatförbund (1)
skal (1/1)
spara (2/2)
frågorfinska (1/1)
kontorstjänster (1/1)
skatteavdrag (1/1)
disk- (1/1)
nybörjare (1/1)
målsättningen (1/1)
inomhus (1/1)
erfarenhetstillägg (1/1)
taget (3/3)
uppstod (1/1)
linkkiRovaniemi (3/3)
beskattning (6/10) Beskattning (4)
tolkningsspråket (1/1)
arbetspensionsutdrag (1/1)
hälsovårdsstiftelses (1/1)
varma (4/4)
bröstsmärtor (1/1)
makas (4/4)
företagsrådgivningen (4/4)
vid (450/450)
ordning (2/2)
biblioteksnätverket (1/1)
psykoterapi (4/4)
var (48/56) Var (8)
bostadsförmedlaren (4/4)
tillfälle (1/1)
människorna (3/3)
barndagvård (8/8)
autonomt (1/1)
arbetsförmåga (1/1)
kandidat- (1/1)
hjärtat (1/1)
parkeringsautomat (1/1)
bestraffning (2/2)
rörelser (1/1)
begäras (2/2)
insjuknar (10/10)
texter (1/1)
innehas (2/2)
intrång (1/1)
idrotts- (1/1)
samjour (1/1)
förmånliga (3/3)
buss (1/1)
kommissionen (1/1)
allmäneuropeiskt (1/1)
utreder (10/10)
vaccineras (1/1)
rättshjälpsbyrå (10/10)
discipliner (1/1)
förvärvsrelaterad (1/1)
åt (22/22)
minst (61/61)
distansundervisning (1/1)
förbereder (3/3)
Kieppi (2/2)
arbetsgivaren (49/49)
Maahanmuuttovirasto (9/9)
torsdagar (2/2)
sjukdomen (1/1)
appen (2/2)
dubbade (1/1)
utveckling (15/18) Utveckling (3)
bastu (6/6)
bekymmer (1/1)
Oy:s (6/6)
undervisningstjänster (2/2)
läggs (1/1)
CV (13/13)
ons. (1/1)
sjukskötarens (2/2)
skolämnen (1/1)
familjfinska (1/1)
händerna (1/1)
undervisningen (26/26)
webbsidor (8/8)
diskriminerat (2/2)
styrkorna (1/1)
nettolönen (1/1)
inte (661/661)
havsvik (1/1)
bostadsägaren (2/2)
föda (3/3)
bastun (4/4)
servicepunkterna (1/1)
operera (1/1)
handelskammare (2/2)
klass (5/5)
varumärkesrätt (1/1)
fattar (15/15)
tillverkningen (1/1)
skaka (1/1)
diskriminerande (2/2)
andelslag (6/6)
egenfinansieringsandel (1/1)
eläke (1/1)
regler (5/5)
förlossningssjukhuset (2/2)
familjemedlem (28/30) Familjemedlem (2)
yrkesinriktade (6/6)
beslutsorganet (1/1)
efternamn (48/48)
ensikoti (1/1)
toimisto.fi (1/1)
serviceproducent (1/1)
centret (5/5)
medlingen (1/1)
ägarbostad (17/20) Ägarbostad (3)
luterilainen (1/1)
notering (1/1)
arbetsuppgiften (4/4)
Europaparlamentsvalet (1/1)
annonser (4/4)
het (1/1)
Konstskolanfinska (1/1)
utrustningen (2/2)
lääkärintodistus (1/1)
riksväg (1/1)
Rooska (1/1)
elevverksamhet (1/1)
slutföra (1/1)
lands (5/5)
äktenskapslagen (1/1)
introduktion (1/1)
arrangerades (1/1)
åtal (1/1)
magistratfinska (1/1)
Korset (6/6)
avsätts (1/1)
arbetslöshetskassorfinska (1/1)
webbplatsfinska (4/4)
uthyrning (1/1)
ID (5/5)
behärskar (2/2)
musikhus (1/1)
oavslutad (1/1)
igen (2/2)
blödningar (3/3)
relationsrådgivningstjänsterfinska (1/1)
invaliditetspension (6/6)
kalkyleras (1/1)
arvsskatt (1/1)
arrangeras (4/4)
öppnad (1/1)
proffs (2/2)
nås (2/2)
medel (17/17)
skilts (1/1)
statsgaranti (2/2)
invandrarens (1/1)
Hedersrelaterat (1/1)
användarråd (1/1)
kartläggningen (14/14)
yrkesutbildade (1/1)
insamlat (2/2)
tatarerna (1/1)
ekonomi- (3/3)
työeläkelaitokset (1/1)
taxitjänster (1/1)
särskilt (15/15)
utbildningslinjer (1/1)
avvecklas (1/1)
hygienen (1/1)
rättigheter (40/41) Rättigheter (1)
visa (12/12)
yrityksen (1/1)
kombineras (1/1)
skiljasfinska (1/1)
verksamhet (40/40)
Kopparbergsvägen (1/1)
Tankkari (1/1)
tittar (1/1)
Schengenstat (1/1)
brottsofferfinska (2/2)
skivor (1/1)
kulturföreningar (2/2)
daghemsdagen (1/1)
förmån (2/2)
tävlingens (3/3)
räkningen (5/5)
Backas (1/1)
specialtjänster (1/1)
enkla (1/1)
asunto (2/2)
hemvårdsstöd (13/13)
Stensvik (1/1)
varningsmärke (1/1)
bondgård (1/1)
persiska (25/25)
territoriet (3/3)
hyrs (9/9)
sommaruniversitetetfinska (1/1)
ortodoxa (13/13)
slovakiska (1/1)
yrkesutbildning (35/36) Yrkesutbildning (1)
Sveriges (2/2)
avgifterna (1/1)
uppföljningen (1/1)
bibliotekets (3/3)
avvisas (1/1)
undersöker (3/3)
nivån (5/5)
estniska (51/51)
Familjeledigheter (1/1)
facket (1/1)
arbetslöshetsförmåner (1/1)
studentkårens (1/1)
regionförvaltningsverk (1/1)
löneutbetalningfinska (1/1)
NA (1/1)
depressionen (1/1)
ungdomsevenemang (1/1)
biljettpriset (1/1)
ungdomsgården (2/3) Ungdomsgården (1)
tolk (40/40)
digital- (1/1)
nätverket (1/1)
kortkurser (1/1)
partiregistret (1/1)
preventionen (1/1)
integreras (1/1)
föräldrars (2/2)
kunskapscentret (1/1)
underhålla (1/1)
brinnande (1/1)
avgiften (4/4)
arbetslivsguide (1/1)
resekort (9/9)
stödja (2/2)
skattedeklarationen (6/6)
finländska (60/64) Finländska (4)
tillståndet (17/17)
resekostnaderna (2/2)
civilståndsintyg (1/1)
efterskott (4/4)
handikappservicen (2/2)
cirka (31/31)
flera (61/61)
tvättstuga (2/2)
miljöområdet (2/2)
samhällslivet (1/1)
sår (1/1)
avsluta (1/1)
skattebyrå (3/3)
kostnadsfri (12/12)
koulutus (3/3)
utfärdas (1/1)
avdragsgill (2/2)
inkräktar (1/1)
kansalaisopisto (2/2)
ungdomsarbetet (3/3)
senast (25/25)
överlåtits (1/1)
könummer (4/4)
handelsplats (1/1)
inträde (3/3)
årstiderna (2/2)
delas (15/15)
helt (5/5)
näringslivet (1/1)
ja (19/19)
Residuum (2/2)
utfärdat (1/1)
Monde (1/1)
vardags- (1/1)
högteknologisk (1/1)
Kejsardömet (1/1)
förbjuda (1/1)
kollektivbostäder (1/1)
mer (418/418)
servicebolag (1/1)
julsånger (1/1)
läkare (35/35)
familjeplanering (5/5)
avdragen (1/1)
stiftas (1/1)
köpeanbud (1/1)
syns (4/4)
boendetjänster (2/2)
nordliga (3/3)
efterfrågan (1/1)
barnfamiljer (7/7)
Sammallahdenmäki (1/1)
hedersrelaterade (2/2)
skattepliktig (2/2)
människovärdet (1/1)
återvända (5/5)
preventivmedel (12/12)
erbjuds (13/13)
Patent- (2/3) patent- (1)
sköts (4/4)
auktoriserad (1/1)
avtalsperioden (1/1)
päivälukio (1/1)
äitiysavustus (2/2)
förskottsuppbördsregistret (2/2)
utgår (3/3)
redogörelse (5/5)
svenskspråkiga (10/10)
grannarna (1/1)
personbeteckning (31/31)
mannens (1/1)
berättar (9/9)
konstnären (1/1)
sorteringen (1/1)
erbjudande (1/1)
byggen (1/1)
bakgaller (1/1)
avlidna (4/4)
veroilmoitus (1/1)
sommarteatern (1/1)
rollen (1/1)
gravt (1/1)
underlättas (1/1)
kontaktinformation (1/1)
fredagar (2/2)
HNS (3/3)
kassakvittot (1/1)
svenskafinska (2/2)
huvudpolisstation (1/1)
jourmottagningfinska (1/1)
föräldramöten (2/2)
offentliggöra (1/1)
medborgare (138/139) Medborgare (1)
lör (1/1)
yrkesutbildningen (1/1)
vårdtillägg (1/1)
brottsligt (1/1)
cykelleder (1/1)
separat (23/23)
yhtiö (1/1)
insjöar (1/1)
nödfall (8/8)
trivsamt (1/1)
anställdafinska (1/1)
starkt (2/2)
ungdomspolitiken (1/1)
utföra (9/9)
gården (1/1)
meta (1/1)
kansalaisuusilmoitus (2/2)
göras (29/29)
vårdnad (16/16)
uppsägningstiden (7/7)
terapibesök (1/1)
problemavfall (1/1)
abonnemang (4/4)
anmälningsblankett (1/1)
märkningen (1/1)
förmåga (2/2)
somaliska (46/46)
civilvigslar (1/1)
fastställs (15/15)
utarbetats (1/1)
halsduk (1/1)
ungas (26/26)
hälsocentralläkarens (1/1)
arbetsgivarförbund (1/1)
bruksvederlag (3/3)
meneefinska (1/1)
strängare (1/1)
systemet (1/1)
stunderna (1/1)
språkkunskaper (27/28) Språkkunskaper (1)
brännskador (1/1)
sjukförsäkringskort (1/1)
kylskåpets (1/1)
åldern (11/11)
liksom (2/2)
Patentti- (1/1)
olja (1/1)
rasistiskt (5/5)
pedagogiska (3/3)
omständigheter (4/4)
utmärkt (1/1)
chatten (2/2)
underhållsbehovet (1/1)
mottagningscentret (1/1)
ersätter (12/12)
Regionförvaltningsverket (2/2)
skyddshemmet (5/5)
flygplats (7/7)
kesäteatterifinska (1/1)
er (8/8)
ll (1/1)
flyttning (1/1)
luopumisilmoitus (1/1)
hälsovårdaren (9/9)
aktiva (5/5)
Sininauha (1/1)
bromsas (1/1)
D (1/1)
pimpelfiske (1/1)
styrker (2/2)
vänskapsförening (1/1)
patients (1/1)
jämställda (3/3)
erityisäitiysraha (1/1)
förlorade (2/2)
meddelar (4/4)
återfå (1/1)
sitter (3/3)
lärokurs (5/5)
skyldigheterna (2/2)
tillställning (1/1)
studierfinska (2/2)
förmögen (1/1)
Chile (1/1)
minimibelopp (1/1)
fakulteterna (1/1)
situationerfinska (1/1)
noga (13/13)
museums (1/1)
företagsservicecentralerna (1/1)
kust (1/1)
barnrådgivningens (1/1)
servicesedlar (1/1)
vårdplats (3/3)
väl (8/8)
anpassningsbara (1/1)
vitsord (5/5)
biologi (1/1)
utför (4/4)
tillfoga (2/2)
immateriella (1/1)
uppstå (1/1)
syn- (1/1)
vårdkostnader (1/1)
polisstationernafinska (1/1)
utsatta (2/2)
yrkesläroanstalter (6/6)
hälsostationsläkare (1/1)
nätbankskoderfinska (1/1)
värmeaggregat (1/1)
befolkningsregistret (5/5)
försvårar (1/1)
hammashoidon (3/3)
tjänstetid (2/2)
stat (4/4)
internet (40/61) Internet (21)
idrottstjänster (5/5)
kunnande (16/16)
fördjupa (1/1)
fritidsverksamhet (1/1)
jympa (1/1)
sjukvårdskort (1/1)
medverka (1/1)
reglerna (4/4)
familjecentret (4/4)
pappersansökan (1/1)
Yrittäjät (1/1)
dagarna (1/1)
smärtjouren (1/1)
allmänhet (10/10)
Päihdelinkki (2/2)
priserfinska (1/1)
ålder (13/13)
vilja (1/1)
aktiv (2/2)
händer (2/2)
informationsmöten (3/3)
motsvarighet (2/2)
svåra (2/2)
samling (1/1)
invånarhusen (1/1)
fatta (5/5)
faderskapserkännande (1/1)
använts (2/2)
blombukett (1/1)
målarfärg (1/1)
kära (1/1)
påbyggnadsnivå (1/1)
grunderna (2/2)
skoldagarna (1/1)
löneperioden (1/1)
flyttfirmorna (1/1)
lägg (2/2)
telefonnumret (2/2)
enda (1/1)
riktad (1/1)
fiska (2/2)
åtagit (1/1)
sköterskan (1/1)
jourmottagningarna (1/1)
övertidstillägg (1/1)
högerextrema (1/1)
dessutom (25/25)
fiskeavfall (1/1)
ämne (3/3)
beskattningsärenden (1/1)
studieprogram (2/2)
kultur- (2/2)
artigt (2/2)
sjukvårdskortet (6/6)
anlänt (2/2)
ställas (3/3)
tandläkare (8/8)
medlemmar (15/15)
motion (26/27) Motion (1)
jourens (1/1)
barnskyddsmyndigheterna (2/2)
barnfinska (7/7)
ockuperade (1/1)
liknande (2/2)
teaterföreställningar (2/2)
nio (5/5)
stämning (1/1)
instanser (2/2)
Förbund (5/5)
indelat (4/4)
mentala (12/12)
närundervisning (1/1)
posta (3/3)
mångkulturella (6/6)
hälsostationsläkaren (1/1)
vattenkannor (1/1)
krisjouren (11/11)
kreditgivningfinska (1/1)
visumärenden (1/1)
utvidgar (1/1)
ungdomsbostadsföreningen (1/1)
utvecklingen (5/5)
sjöfästning (1/1)
föddes (1/1)
anhålla (1/1)
läroplanen (1/1)
psykiska (6/6)
Vantaa (1/1)
arbetssätt (1/1)
välartat (1/1)
innebära (1/1)
anledning (5/5)
bistånd (1/1)
sjukvårdstjänster (5/5)
försäljningsställen (1/1)
utan (101/101)
maka (31/31)
insjuknat (1/1)
sida (270/270)
registrerat (12/12)
misstänka (1/1)
dansa (3/3)
ledamöter (5/5)
handläggningsavgift (1/1)
grader (3/3)
patientombudsmannen (2/2)
51:a (2/2)
vräka (1/1)
personalen (5/5)
demensfinska (1/1)
berättelse (1/1)
tingsrättenfinska (1/1)
affärsresa (1/1)
godtas (1/1)
Kilo (2/2)
myndighetsärenden (1/1)
sökte (1/1)
annans (2/2)
trafikfinska (1/1)
medborgarskapfinska (3/3)
bruksvederlaget (2/2)
kommunernafinska (2/2)
utrustning (3/3)
säkerhetsanvisningar (1/1)
jobbannonsen (3/3)
strävar (3/3)
Ilmonet.fi (1/1)
genetiska (1/1)
tänka (2/2)
aktivt (4/4)
fjärde (13/13)
liten (11/11)
arbetslöshetsförmånen (2/2)
arbetsmiljö (1/1)
omfatta (5/5)
bouppteckningen (3/3)
fast (10/10)
servicepunkter (1/1)
land (140/140)
förhandlare (1/1)
åtgärdande (1/1)
stället (2/2)
veronpalautus (2/2)
-trivsel (1/1)
byggherren (1/1)
skattar (1/1)
färdtjänster (1/1)
språkkurser (3/3)
ungdomarfinska (2/2)
varan (1/1)
responsen (1/1)
integrationsspråk (1/1)
dödsfallet (1/1)
bevilja (1/1)
RFV (1/1)
hänt (1/1)
kollektiv (1/1)
starka (2/2)
finansieringen (4/4)
lekparksträffar (1/1)
brottsoffrets (1/1)
HelMet (3/4) Helmet (1)
uppbära (1/1)
Mårtensdal (1/1)
rösta (16/16)
tidsbokningssystem (1/1)
isen (7/7)
födas (1/1)
R3 (2/2)
studentskrivningarna (1/1)
stödjer (5/5)
kärren (1/1)
kontaktar (3/3)
förskoleundervisningfinska (3/3)
högt (4/4)
timmar (14/14)
taket (1/1)
fastlagen (1/1)
ammattikorkeakoulu (4/4)
livet (11/12) Livet (1)
rehabilitering (42/43) Rehabilitering (1)
brottsanmälanfinska (1/1)
lära (21/21)
olydiga (1/1)
skogsindustrin (1/1)
alternativt (2/2)
varifrån (1/1)
räntestödetfinska (1/1)
arbetskollektivavtal (1/1)
skolläkaren (3/3)
äktenskapslagenfinska (1/1)
studiestöd (8/8)
sökandena (1/1)
förhållandena (1/1)
lånetiden (1/1)
Östersjön (1/1)
köp (5/5)
miljö- (1/1)
väder (1/1)
affärsidé (1/1)
parrådgivning (1/1)
specialfinansieringsbolag (1/1)
universitetsexamen (2/2)
deltagarna (1/1)
Sodankylä (1/1)
anställningsskyddet (1/1)
fackförbundsverksamhetfinska (2/2)
spårvagnarna (1/1)
praktiken (5/5)
liikenne (1/1)
klient (1/1)
European (1/1)
skolresestödetfinska (1/1)
tidningar (9/9)
jaktfinska (1/1)
webbsida (2/2)
döma (1/1)
arbetsuppgifterna (2/2)
arbetspension (6/6)
mervärdesskatt (3/3)
skulle (9/9)
stadgas (3/3)
utvecklingsstörning (1/2) Utvecklingsstörning (1)
litauiska (1/1)
skattenumret (3/3)
öppen (13/13)
mycket (66/66)
julskinka (1/1)
tystnadsplikt (2/2)
anslutning (8/8)
individuell (1/1)
anhörigas (1/1)
närståendevård (6/6)
trauma (1/1)
vanliga (12/12)
överskridits (1/1)
klubben (2/2)
cykel (1/1)
anlitar (1/1)
regionen (3/3)
ehkäisyneuvonta (1/1)
specialundervisning (5/5)
avläggs (1/1)
pensionens (1/1)
länsbaserade (1/1)
förebyggandet (1/1)
bidragens (1/1)
dagstidningar (2/2)
verka (2/2)
utomlands (61/61)
oljud (3/3)
syskon (4/4)
förskola (2/2)
Schengenländerna (1/1)
vaccinerar (1/1)
universitetskurser (1/1)
beskattningsbara (3/3)
ingåtts (5/5)
körkortfinska (1/1)
källa (1/1)
bygget (1/1)
biografer (3/3)
samarbetsmöjligheter (1/1)
bedömningen (1/1)
Osviitta (1/1)
Unescos (1/1)
frånvaron (1/1)
skyddshus (10/10)
reparera (1/1)
påbörjas (2/2)
medlemsfamiljerna (1/1)
hundratals (1/1)
månaders (5/5)
ledda (2/2)
bilskatten (1/1)
ombyggnadsarbeten (1/1)
vetenskap (1/1)
källan (1/1)
sång (1/1)
häradsskrivare (1/1)
fyllda (1/1)
rimligt (2/2)
bolaget (1/1)
framställning (1/1)
verokortti (3/3)
obetalda (2/2)
Miehen (6/6)
bokat (4/4)
hyresgaranti (1/1)
YH (2/2)
kräva (10/10)
älvarna (1/1)
hektar (1/1)
Estland (1/1)
mörkare (1/1)
Kipinä (2/2)
gymnasiet (21/21)
cykeln (1/1)
formulerad (1/1)
kl (73/73)
servicepunkten (3/3)
tvingar (1/1)
skattmyndigheten (1/1)
antibiotika (1/1)
utbytesstudier (1/1)
unionen (6/6)
ordkonst (1/1)
tillsvidareanställning (1/1)
osakeyhtiö (1/1)
representerar (6/6)
skaffat (1/1)
Vandafinska (1/1)
grundade (2/2)
tietopankki (1/1)
prick (1/1)
faderskapspenning (3/3)
egna (44/44)
työterveyshuolto (1/1)
förälder (36/36)
språkexamina (5/5)
nuorisoasema (1/1)
försätts (1/1)
ber (1/1)
ärvs (1/1)
bostadsrättsavgifter (1/1)
webbankkoderna (1/1)
avslås (1/1)
bindestreck (1/1)
arrangerar (1/1)
kommunerer (1/1)
dagvårdsplats (8/8)
girering (1/1)
styrka (9/9)
IHH (1/1)
kallas (12/12)
Esbobor (1/1)
skiftesvård (1/1)
planerad (1/1)
riksdagsledamot (1/1)
vigsel (11/11)
träffarna (1/1)
finskspråkigt (2/2)
patientjournalen (1/1)
kör (1/1)
arbetspensionsförsäkringarna (1/1)
varit (22/22)
öka (2/2)
flyttanmälan (3/3)
entrédörren (2/2)
överföringen (1/1)
urologisk (1/1)
betalningar (3/3)
klinikstiftelsens (2/2)
produktionsmedel (2/2)
slotten (2/2)
intresserade (6/6)
etniskt (7/7)
hyvinvoinnin (1/1)
nuortenkeskus (2/2)
koulupsykologit (1/1)
landet (32/32)
lärokursen (2/2)
skötare (5/5)
preliminär (1/1)
påföljder (1/1)
B2 (1/1)
biträdande (1/1)
ungdomsgårdar (5/5)
respektive (2/2)
organisationen (1/1)
www.infopankki.fi (1/1)
receptet (1/1)
statsförvaltningens (5/5)
hantera (2/2)
hälsostationer (10/10)
invandrarmänfinska (1/1)
tas (23/23)
stadiluotsi (1/1)
gynekolog (4/4)
föremål (2/2)
trafikeras (1/1)
tillfrisknande (1/1)
museerna (4/4)
Varia (3/3)
anlita (14/14)
räkningar (2/2)
eläkevakuutus (2/2)
gård (1/1)
Rovanapa (2/2)
svarat (1/1)
skadar (1/1)
stiftelsens (2/2)
konstundervisningfinska (1/1)
servicehus (5/5)
yrkesstudier (1/1)
mobilabonnemang (1/1)
giltiga (2/2)
barnpassning (1/1)
måste (206/206)
förra (1/1)
räknar (1/1)
föreningarfinska (1/1)
styrelsemedlem (1/1)
vårdinrättning (2/2)
underhåller (1/1)
meddelats (1/1)
begäran (6/6)
tempus (1/1)
hindersprövningen (6/6)
förrättas (14/14)
grupps (1/1)
uppförandet (1/1)
ungdomsväsendet (1/1)
lagarna (5/5)
synnerhet (1/1)
fritidsintressen (3/3)
staterna (1/1)
rötterna (1/1)
ingrepp (1/1)
könsminoriteterfinska (1/1)
aning (1/1)
stads (61/61)
webbankkoder (4/4)
metallindustrin (1/1)
läsår (4/4)
Creative (1/1)
sökmotorns (2/2)
kvotflyktingar (8/8)
adopterar (1/1)
Västerkulla (1/1)
Sovjetunionens (1/1)
tolktjänst (2/2)
erfarenhet (2/2)
arbetslivets (1/1)
bevåg (1/1)
stadsdirektören (1/1)
passar (7/7)
samtalar (3/3)
medlemsländer (1/1)
presenteras (3/3)
motsätter (2/2)
pratar (4/4)
längre (23/23)
internettjänsten (1/1)
Kluuvi (1/1)
staten (8/8)
korta (4/4)
original (6/6)
tunnustaminen (1/1)
avgjorts (1/1)
reservationsavgifter (1/1)
agerar (1/1)
utbildade (4/4)
prepositioner (1/1)
samfundet (1/1)
parkeringsbiljett (1/1)
dagpenningens (1/1)
advokatförbundfinska (1/1)
fara (6/6)
lagringsavgifter (1/1)
ägt (1/1)
hobbymöjligheter (2/2)
Företagsfinlands (2/3) FöretagsFinlands (1)
dör (6/6)
terapi (2/2)
sex (22/22)
elevernas (3/3)
betalningsdagar (1/1)
sjukdomstid (2/2)
närvarar (1/1)
visering (1/1)
tacka (2/2)
bereds (1/1)
yrkesexamenfinska (1/1)
nationell (1/1)
lagrar (1/1)
juristen (1/1)
tandvårdens (2/2)
anmälningsdagen (2/2)
dricks (1/1)
minimikraven (1/1)
ovanlig (1/1)
dennes (4/4)
lantdagsmannen (1/1)
respektera (1/1)
hyresdeposition (2/2)
bemötande (3/3)
Rex (2/2)
områden (17/17)
privata (45/45)
ursprung (12/12)
juristhjälp (1/1)
tyngdpunkt (1/1)
tfn (16/17) Tfn (1)
register (1/1)
tvinga (8/8)
arbetsinkomst (2/2)
årervinns (1/1)
resor (2/2)
dubbelexamen (1/1)
formella (1/1)
bostadsförmedlingen (1/1)
hyran (14/14)
beslutsfattarna (1/1)
specialutbildning (1/1)
bland (38/38)
fortsättningskriget (1/1)
delen (10/10)
resten (3/3)
bästa (11/11)
bekräftande (1/1)
receptfinska (1/1)
fönstret (1/1)
bostadssökande (1/1)
utbildningsväsendetfinska (1/1)
Helsinkis (1/1)
halvt (1/1)
l (3/3)
rehabiliteringsinrättning (1/1)
hautaustoimisto (2/2)
text (1/1)
våren (14/14)
elektronisk (5/5)
fullständigt (1/1)
hälsocentralsjouren (1/1)
verkliga (2/2)
tillståndstjänstenfinska (1/1)
biljetter (2/2)
utses (3/3)
resekorten (1/1)
CD- (1/1)
läst (4/4)
hindersprövning (5/5)
gjort (5/5)
avgiftsfria (8/8)
pappersformat (1/1)
översättas (3/3)
provar (1/1)
organisationer (15/15)
via (103/103)
samman (2/2)
närskolan (2/2)
Nuorisosäätiö (2/2)
laddat (1/1)
rådgivningsställe (1/1)
hälsostationen (38/38)
kommunsidorna (1/1)
elbolags (1/1)
Klimatet (1/2) klimatet (1)
grammatikövningar (1/1)
skatt (21/21)
punktskriftsböcker (1/1)
storlek (16/16)
takt (2/2)
namnlag (1/1)
asunnotfinska (1/1)
problem (83/90) Problem (7)
Kansa (1/1)
hälscentralsavgifter (1/1)
binder (2/2)
återhämtningen (3/3)
universitet (43/48) Universitet (5)
kouluterveydenhoitaja (1/1)
industristad (1/1)
omhändertagande (1/1)
fordon (1/1)
mylla (1/1)
migration (1/1)
skräpa (1/1)
YTHS (1/1)
Insurance (1/1)
engelskspråkig (6/6)
gick (2/2)
utrikespolitiken (1/1)
person (64/64)
Vuokra (1/1)
Norge (7/7)
tolken (13/13)
rusmedel (2/2)
hindrar (1/1)
legaliserad (2/2)
säkerhetstjänster (1/1)
barnrådgivningsbyråns (1/1)
mängd (5/5)
metodstudier (2/2)
Alkoholister (2/3) alkoholister (1)
värdesätts (4/4)
utsätta (1/1)
baserade (1/1)
vakuutusyhtiö (1/1)
sjukvårdstjänsterna (4/4)
uppsägningsvillkor (3/3)
genomsnitt (4/4)
gravid (7/7)
löneintyg (4/4)
Kotoutumiskeskus (1/1)
baltiska (1/1)
sommaruniversitetet (2/2)
säkerställer (1/1)
lokalerna (1/1)
kommuner (20/20)
servicebostadsgrupp (1/1)
småbarnspedagogik (11/11)
halt (2/2)
sak (5/5)
lägenheter (1/1)
bolagsavtal (1/1)
tjänsteleverantör (1/1)
misslyckades (1/1)
studieregisterutdrag (1/1)
behöver (266/270) Behöver (4)
bifogas (1/1)
boendeträffpunkter (1/1)
socialskyddsavtal (2/2)
framför (1/1)
barnrådgivningsbyrån (1/1)
bortgång (1/1)
förvärvsarbetande (1/1)
Sveaborgs (1/1)
skogar (1/1)
utarbetas (5/5)
hyresdepositionen (3/3)
firandet (1/1)
lapsettomuusklinikka (1/1)
sund (1/1)
självstyre (2/2)
fritidsaktiviteter (3/3)
grundskolebaserad (4/4)
Kvarkens (1/1)
Stadin (4/4)
energibesparingslampor (1/1)
familjecenter (1/1)
skriven (1/1)
vidtar (1/1)
akut (22/22)
misstänkt (1/1)
tidiga (3/3)
läroämnen (4/4)
ammatti- (3/3)
yrkesval (1/1)
upphovsmannen (1/1)
sälja (6/6)
studeranden (7/7)
skräp (1/1)
skilsmässa (50/54) Skilsmässa (4)
förbättra (12/12)
magisterprogram (4/4)
misstanken (1/1)
hemifrån (2/2)
ihåg (25/25)
steril (2/2)
bygg (1/1)
undervisningenfinska (2/2)
franskan (1/1)
rådgivningstjänsten (1/1)
observera (3/3)
ramper (1/1)
normala (1/1)
vistats (6/6)
flyttsakerna (1/1)
Metropolias (1/1)
patienter (1/1)
religionssamfunds (2/2)
Abfinska (1/1)
Uusi (1/1)
vuxengymnasiet (5/5)
piller (2/2)
Helsingfors (169/169)
utbyten (1/1)
Suomen (12/13) suomen (1)
gamla (8/9) Gamla (1)
nyttiga (2/2)
välsignas (1/1)
roll (2/2)
SOS (1/1)
färdtjänsten (1/1)
läkarstationer (4/4)
EVK (1/1)
kreditkort (3/3)
bl.a. (7/7)
skrivfärdigheter (1/1)
undersökning (8/8)
anmälas (5/5)
mousserande (1/1)
samma (72/72)
institutioner (2/2)
Karleby (56/56)
vars (20/20)
språken (5/5)
könsminoriteters (1/1)
ska (417/417)
ordningsreglerna (7/7)
sköter (23/23)
kränkande (1/1)
Easyfinnishfinska (1/1)
besöksförbud (3/3)
riktnummer (1/1)
grundskolans (12/12)
sairauspäiväraha (2/2)
viktigaste (9/9)
minoritetsspråk (1/1)
anknyter (4/4)
rättsskyddsförsäkring (1/1)
van (1/1)
hemfriden (1/1)
bussbiljetter (1/1)
undervisningstillstånd (1/1)
eduskunta (2/2)
samverkan (1/1)
diskmaskin (1/1)
lönespecifikationen (2/2)
Suomenlinna (1/1)
sjukledigheten (3/3)
skyldigheter (23/23)
personbeteckningen (7/7)
apotekens (1/1)
dömer (1/1)
abortti (1/1)
läckaget (1/1)
privatskolor (1/1)
batterier (1/1)
fuktisolering (1/1)
betjäning (3/3)
VAU (1/1)
reseersättning (1/1)
utbildningsväsendet (2/2)
hälsovårdsministeriets (3/3)
svårt (17/17)
förebyggande (6/6)
hälsovårdscentralen (7/7)
handarbete (4/4)
stöda (4/4)
parets (1/1)
närståendevårdare (1/1)
tävlingsarrangören (1/1)
skolornas (2/2)
läroavtal (3/3)
lätta (1/1)
avgiftsbelagt (4/4)
regionkontor (1/1)
undgås (1/1)
löntagare (1/1)
kärnkompetens (2/2)
efterlevandes (1/1)
måltidsstöd (1/1)
boendekostnaderna (6/6)
tidigt (6/6)
förblir (3/3)
berusad (1/1)
tideräkningen (1/1)
ladda (7/7)
vardagkvällar (1/1)
delgivits (1/1)
pimpla (2/2)
fastighetsägare (1/1)
måltider (4/4)
betjäna (1/1)
startas (1/1)
folkomröstningar (1/1)
resesättet (1/1)
arbetssökande (25/25)
hälsocentral (1/1)
mallarfinska (1/1)
toimipiste (1/1)
lördagar (1/1)
fyllde (1/1)
moderskapspenningperiodens (1/1)
får (399/399)
din (511/511)
inträffat (2/2)
anvisning (1/1)
frysen (1/1)
följd (5/5)
finskspråkig (3/3)
sittunderlag (1/1)
kuntoutuslaitos (1/1)
klicka (1/1)
vädret (2/2)
upphöra (2/2)
allemansrätten (2/2)
pensionfinska (1/1)
förvaltningsdomstolen (5/5)
moderskapsledighet (2/2)
beskattningen (24/24)
Näringsliv (3/3)
förmedling (1/1)
livmoderhalscancer (2/2)
rasistiska (2/2)
yttra (1/1)
rf (11/11)
skaffas (1/1)
islamska (1/1)
kommanditbolag (4/4)
sjukhusjouren (1/1)
seurakunnan (1/1)
Päivystysapu (1/1)
hemkommunen (3/3)
föreningsverksamhet (2/2)
anhörigvård (1/1)
yta (1/1)
påverkat (1/1)
vanligen (46/46)
annorlunda (2/2)
domstolen (4/4)
kielenä (1/1)
Vionoja (1/1)
hyresvärdar (5/5)
allmäneuropeisk (1/1)
påverkas (7/7)
berättigar (2/2)
musikverksamhet (1/1)
fem (24/24)
identitet (14/14)
tonåringar (1/1)
motsvarande (5/5)
yrkesutbildningar (1/1)
samboförhållandet (6/6)
myndig (5/5)
självständighetsdagen (1/1)
Lappland (6/6)
bolagsordningen (1/1)
utomstående (3/3)
tobak (1/1)
uppstår (5/5)
bilskatt (1/1)
intressanta (1/1)
hyressed (1/1)
tjänsteprocesserna (1/1)
bekantskaper (1/1)
klär (1/1)
löneanspråk (1/1)
ugriska (1/1)
kustregionerna (1/1)
bröstcancer (2/2)
ändring (1/1)
TyEL (1/1)
ämnar (2/2)
kondylom (1/1)
vårdbidrag (1/1)
studiemöjligheter (5/5)
MB (10/10)
uppleva (1/1)
ståt (1/1)
återvändandefinska (1/1)
hörsel (2/2)
abonnemanget (1/1)
betalningsanmärkning (2/2)
kommandiittiyhtiö (1/1)
nödnumretfinska (1/1)
plastkasse (2/2)
vardagen (7/7)
ry. (1/1)
skatter (9/9)
gifta (23/23)
fött (3/3)
parternas (1/1)
avancerad (1/1)
vågar (2/2)
mening (1/1)
familjeförening (2/2)
vinster (1/1)
sysselsättningsstöd (2/2)
barnförhöjningen (1/1)
utformas (1/1)
krisjour (3/3)
visning (1/1)
riksdagsledamöter (1/1)
yrken (11/11)
sökt (3/3)
garantipensionens (1/1)
tung (1/1)
tillfälligt (21/22) Tillfälligt (1)
museet (3/3)
stödspråkfinska (1/1)
demokratiska (1/1)
ungdomarna (2/2)
svara (1/1)
kontaktade (1/1)
löptid (1/1)
fest (3/3)
-Förbundet (1/1)
rädda (1/1)
landsbygd (1/1)
ibland (11/11)
bostaden (62/62)
bankonto (1/1)
skatteåterbäring (4/4)
lågkonjunkturen (1/1)
bestå (6/6)
vandrarhem (1/1)
samtliga (11/11)
trafik- (1/1)
beter (2/2)
behovsprövat (2/2)
reliefbilder (1/1)
använda (79/79)
mödra- (8/8)
graviditet (10/10)
serviceboendet (2/2)
Studentkårers (1/1)
yksityisen (1/1)
läkarcentral (1/1)
sättas (1/1)
studieplatsen (1/1)
finländskt (5/5)
hobbyverksamhet (5/5)
Europaparlamentsval (4/4)
definierar (1/1)
fre (22/22)
endera (4/4)
personerlinkkiEsbo (1/1)
skidåkning (2/2)
förlossningssjukhus (1/1)
webbenkäter (1/1)
köpare (2/2)
tidskrifter (3/3)
Luksia (1/1)
betalningstiden (3/3)
släckningsfilt (2/2)
hälsovårdstjänster (23/26) Hälsovårdstjänster (3)
beviljandet (1/1)
bort (4/4)
linkkiLapplands (1/1)
kaffesump (1/1)
EMMA (1/1)
måltidservice (1/1)
center (5/5)
försämrar (1/1)
växter (1/1)
flyttrörelsen (1/1)
fax (3/3)
yrkena (1/1)
toimisto (4/4)
hälsotillstånd (7/7)
oppilaitos (1/1)
antalet (5/5)
vinterskor (1/1)
ned (6/6)
huvudhälsostation (1/1)
familjeterapi (1/1)
kvalifikationer (4/4)
affärsidén (2/2)
Flerspråkiga (2/2)
expert (1/1)
grannkommunen (1/1)
öst (2/2)
rusmedelsberoendefinska (2/2)
Pulkamontiefinska (1/1)
informationsservice (1/1)
bosättningsland (1/1)
hobbyklubbar (1/1)
beträda (2/2)
yrkesvägledning (1/1)
mån. (1/1)
hemspråksundervisning (5/5)
året (19/19)
MIELI (2/2)
köpta (1/1)
föräldralediga (1/1)
representeras (1/1)
gå (36/36)
personal (2/2)
teaterstad (1/1)
behöva (6/6)
abort (8/9) Abort (1)
larm (1/1)
problematiska (5/6) Problematiska (1)
Wilma (6/6)
musikgrupper (1/1)
hurdana (6/6)
gör (30/30)
skolväsendet (1/1)
kontakter (2/2)
förändring (1/1)
verotoimisto (3/3)
yrkesbenämning (1/1)
vistelse (9/9)
musikskolor (1/1)
rödbetssallad (1/1)
utvecklingsstadium (1/1)
allmän (8/9) Allmän (1)
faktorer (2/2)
telefontid (1/1)
saken (9/9)
besluta (10/10)
kontrollen (1/1)
dess (18/18)
tempel (1/1)
kollektivtrafikens (5/5)
Kemi (1/2) kemi (1)
avtalade (2/2)
ung (7/7)
organisationsverksamhet (1/1)
språkversioner (1/1)
Livsmedelsverket (1/1)
inriktningar (1/1)
realiseringen (1/1)
festivalen (1/1)
demokratin (1/1)
narkomaanit (1/1)
uppvärmningen (1/1)
hobbyer (4/4)
utlänningarengelska (1/1)
tolkning (3/3)
familjemedlems (1/1)
slogs (1/1)
försörjningsförutsättningen (2/2)
Bottniska (2/2)
vigselfinska (2/2)
psykologhjälp (1/1)
trädgårdsskötsel (1/1)
tillståndsenhet (1/1)
spela (4/4)
sker (14/14)
verksamhetsställen (9/9)
jobba (2/2)
tätorter (2/2)
sammanhängande (1/1)
www.kopiosto.fi (1/1)
rajoitetusti (1/1)
kaffepaus (2/2)
trähus (1/1)
arbetarskydd (2/3) Arbetarskydd (1)
skydda (3/3)
bestämmelser (2/2)
omskurits (2/2)
delar (11/11)
statsborgen (1/1)
förbrukning (3/3)
överklagande (1/1)
handlingen (2/2)
grenar (3/3)
brutit (2/2)
ministrarna (1/1)
uppsägningen (1/1)
förutsättningarna (3/3)
undersökningen (3/3)
kompletterande (2/2)
behandlas (28/28)
första (40/40)
betydande (1/1)
startpeng (5/5)
tidskriften (1/1)
universitets (3/3)
hemvården (2/2)
gälla (2/2)
motivera (1/1)
flyttade (6/6)
Kannus (1/1)
arbetsgivarens (4/6) Arbetsgivarens (2)
vuxnafinska (3/3)
ringa (58/58)
varierar (18/18)
hälsostation (37/37)
alkuomavastuu (1/1)
lokal- (1/1)
lever (4/4)
planerar (10/10)
jourtidsbeställning (1/1)
kremeras (1/1)
valts (1/1)
föräldrapenningsperioden (1/1)
gripa (1/1)
HRT:s (2/2)
emellan (1/1)
tolkningstjänsten (1/1)
Nupoli (4/4)
organiserade (1/1)
esteiden (3/3)
jakt (2/2)
mataffären (1/1)
hudfärg (3/3)
arbetslöshetsförmånfinska (1/1)
viktigast (1/1)
yrkesinstitut (8/8)
försäkring (7/7)
företagshälsovård (8/9) Företagshälsovård (1)
kämpades (1/1)
krisområden (1/1)
förmögnare (1/1)
ännu (10/10)
ramen (1/1)
förödmjukande (1/1)
ungdomstjänsterfinska (1/1)
återvinningsstationer (1/1)
förväg (22/22)
fiskeredskap (1/1)
bevisas (4/4)
turvatalo (3/3)
hallinto (1/1)
egendomsfördelning (1/1)
universitetsstudier (3/3)
psykoterapitjänst (1/1)
skolhälsovårdarna (1/1)
Renlunds (1/1)
omsorgsfullt (2/2)
varhaiskasvatuspäällikkö (1/1)
underskridas (1/1)
viktiga (7/9) Viktiga (2)
norr (1/1)
inlärning (4/4)
samtalspriset (1/1)
skydd (12/12)
högljudd (1/1)
km (1/1)
betydelse (1/1)
insatt (2/2)
påvisas (1/1)
besvaras (2/2)
fortare (1/1)
anledningar (1/1)
fordonsskatten (1/1)
TE (73/74) te (1)
först (50/50)
bosatta (16/16)
fostrets (2/2)
Pejas (2/2)
kommuntilläggfinska (1/1)
utländsk (15/16) Utländsk (1)
uppgifterna (12/12)
befolkningsdatasystem (4/4)
uppdragsavtal (2/2)
tala (14/14)
friluftsmuseumfinska (1/1)
användarna (4/4)
åligger (2/2)
kärnkraftverket (3/3)
smittats (1/1)
tilltalar (1/1)
därmed (2/2)
begära (14/14)
resmålen (1/1)
längs (1/1)
inkomstrelaterad (9/9)
transporttjänst (1/1)
arvodet (1/1)
stranden (1/1)
näringsbyråerna (4/4)
tandborstar (2/2)
tjänstemannafinska (1/1)
lagstadgade (1/1)
is (1/1)
ytterligare (9/9)
oikeudet (1/1)
arbetstid (10/10)
sopsorterar (1/1)
Begravningbyråers (1/1)
landfinska (1/1)
arbetslivet (20/20)
överenskommits (3/3)
vem (15/15)
högklassiga (1/1)
institution (1/1)
sähköinen (1/1)
trafik (3/3)
ansökningsblankett (9/9)
uhrien (1/1)
möjligt (41/41)
socialtjänsterna (2/2)
erhållit (2/2)
bedriva (1/1)
hundra (1/1)
kondomer (1/1)
innehåller (14/14)
Alexandersgatan (1/1)
cirkuskonst (2/2)
årligen (1/1)
utskrivna (1/1)
förklarade (1/1)
italienska (15/15)
mångsidiga (3/3)
regeringen (2/2)
utgift (1/1)
nationalmuseumfinska (1/1)
ytan (1/1)
löner (2/2)
konstaktiviteter (1/1)
gått (10/10)
livförsäkring (1/1)
anställda (45/45)
Aalto (2/2)
läger (3/3)
hobbygrupper (1/1)
musiker (1/1)
aldrig (2/2)
operation (2/2)
lämplighet (1/1)
utbytesstudent (2/2)
Schengenvisum (1/1)
läkarstation (14/14)
stationen (1/1)
livlig (1/1)
tillhör (11/11)
tukiverkko (1/1)
betalning (1/1)
huvudjärnvägsstation (1/1)
Schweiz (31/31)
Dublinprocessen (1/1)
förenings (1/1)
skolhälsovården (2/2)
anställningen (9/9)
begär (2/2)
infopankki (1/1)
område (28/28)
del (65/65)
motionfinska (1/1)
hänvisas (1/1)
utdrag (3/3)
Finavia (1/1)
erillinen (1/1)
organisation (4/4)
avancerade (1/1)
vaccinationerna (2/2)
tvärtom (1/1)
hemvårdsavgiften (1/1)
HIV (2/2)
sjukdomsattack (1/1)
Apostilleintyg (1/1)
heminkvartering (1/1)
pensionärsrabatten (1/1)
bilda (1/1)
verksamhetsstället (1/1)
kulturhistoria (2/2)
fungerar (5/5)
nättjänsterna (2/2)
Banvägen (1/1)
drogs (1/1)
förnamn (1/1)
identitetshandling (6/6)
Åbo (7/7)
häxor (1/1)
resurscenter (1/1)
krigsskadeståndet (1/1)
kvälls- (2/2)
mitt (9/9)
grekiska (2/2)
länkar (5/5)
socialservice (1/1)
affärsförhandlingar (1/1)
förslag (3/3)
samfundfinska (2/2)
uppgift (8/8)
tisdag (1/1)
vice (1/1)
minimilönerna (1/1)
barn (315/319) Barn (4)
diskuterar (2/2)
naturcenter (1/1)
nivå (7/7)
fackevenemang (1/1)
hemsjukvård (1/1)
utbildningsanordnare (1/1)
regnbågsfamiljerfinska (1/1)
syssla (2/2)
CV:t (2/2)
påsken (1/1)
olycksfallsstation (2/2)
tv (5/6) TV (1)
vintern (7/7)
ersättningsgill (1/1)
työsuojelun (1/1)
upprepa (1/1)
flerfaldigt (5/5)
understöds (1/1)
yrkeshögskola (18/18)
fortbildning (5/5)
fars (1/1)
igång (2/2)
vinterkriget (1/1)
andras (3/3)
diskrimineringsombudsmannens (2/2)
terapin (2/2)
Haartmanska (4/4)
beviljades (3/3)
Finlandfinska (28/28)
Korsets (1/1)
föreningsmöten (1/1)
tjänsteleverantörers (1/1)
skattefria (1/1)
friare (1/1)
finländarna (19/19)
utom (4/4)
köpas (6/6)
rutter (5/5)
strid (1/1)
Böle (4/4)
kvinnorna (3/3)
minskar (3/3)
uppdrag (3/3)
stödpersonen (1/1)
bruk (3/3)
amorteras (1/1)
stadens (53/53)
hyresvärdarnas (1/1)
arkivet (1/1)
försäkringsbolaget (1/1)
ansvariga (5/5)
föräldradagpenning (5/5)
inledande (27/27)
detalj (1/1)
läggning (6/6)
socialskyddet (3/3)
näringstjänsten (1/1)
lekparker (3/3)
Ullava (3/3)
hälsorelaterade (1/1)
initiativtagande (1/1)
hobby (7/7)
samboskap (1/1)
tandvård (19/19)
finansieringsbolag (1/1)
svalt (2/2)
perheneuvonta (1/1)
hyötyliikunta (1/1)
hörseln (1/1)
guld (1/1)
opetuksen (1/1)
aktuell (4/4)
daghemsföreståndarna (2/2)
miljoner (1/1)
sydkusten (1/1)
utlänningsbyrån (3/3)
nettopalkka (1/1)
transvestiter (1/1)
missbrukstjänster (1/1)
Inre (4/4)
lägenhetshotell (2/2)
konstarter (3/3)
Hautaustoimistojen (1/1)
toiminimi (2/2)
stulits (1/1)
förbudet (1/1)
exempel (355/355)
ungdomsverksamheten (1/1)
PISA (1/1)
kallare (1/1)
dit (6/6)
innan (75/75)
system (3/3)
opintolinja (1/1)
kvarskatt (3/3)
måltidstjänster (1/1)
franska (60/60)
sålt (1/1)
priser (5/5)
grundskoleinstitutionen (1/1)
hens (1/1)
värme (1/1)
socialhandledningfinska (1/1)
medborgares (7/7)
flyttsaker (4/4)
innehållen (1/1)
separation (1/1)
työkyvyttömyyseläke (1/1)
mielenterveysseuran (1/1)
koulu (2/2)
alkoholdrycker (2/2)
inreseförbud (2/2)
duger (3/3)
fre. (1/1)
bestäms (6/6)
taasengelska (1/1)
kontaktspråk (1/1)
institut (6/6)
mödrahemsverksamheten (1/1)
postadress (1/1)
familjsvenska (1/1)
examensnivå (1/1)
rehabiliteringsbeslut (1/1)
bussbolag (1/1)
rökfria (1/1)
fotografi (1/1)
Väestörekisterikeskus (1/1)
kvalitet (2/2)
arbetets (2/2)
examensstuderande (2/2)
Herman (1/1)
beredd (1/1)
järnaffärer (1/1)
boendetfinska (1/1)
kompletterar (2/2)
Esbos (1/1)
jämställdhetsnämnden (4/4)
äventyra (1/1)
Vandatillägget (1/1)
kuntoutus (2/2)
allra (2/2)
avlidne (4/4)
skärgårdenfinska (1/1)
oväntat (2/2)
köparen (2/2)
medeltiden (1/1)
mån (16/16)
milda (1/1)
kurs (4/4)
uppehållstillstånden (1/1)
sorts (2/2)
lovat (2/2)
behandlar (4/4)
koncentrationssvårigheter (1/1)
bärbar (1/1)
resehandling (2/2)
varuhus (1/1)
erhålla (3/3)
återkallar (2/2)
annonsen (2/2)
bedrivit (1/1)
bostadslösafinska (2/2)
reparation (1/1)
utvisad (1/1)
sen (1/1)
kotihoito (1/1)
demonstration (1/1)
träd (3/3)
eventuella (7/7)
hälsocentraler (1/1)
genus (1/1)
grannmedlingfinska (1/1)
lääkäri (2/2)
kvotflykting (4/4)
dokument (4/4)
finansiärerna (1/1)
kastrullock (1/1)
Smith (2/2)
tillväxtföretagare (2/2)
äktenskapshinder (6/6)
rådgivningstjänsterna (3/3)
ämnena (1/1)
utomlandsfinska (2/2)
andraspråk (3/3)
festmat (1/1)
avsnittet (1/1)
tyska (38/38)
eija.kyllonen (1/1)
lånesumman (1/1)
yrkesinstitutet (1/1)
frågorna (1/1)
upplösning (2/2)
äänioikeusrekisteri (1/1)
sambon (4/4)
Kriscentret (1/2) kriscentret (1)
metrostationer (1/1)
beräkna (3/3)
invånarlokalen (1/1)
ventilation (1/1)
överskrids (1/1)
skyddshusfinska (2/2)
Business (5/5)
patienten (4/4)
ämbetsbevis (2/2)
personers (3/3)
slutade (1/1)
sökandes (1/1)
ansvarar (12/12)
lite (11/11)
nödvändig (3/3)
födelseattest (6/6)
sosiaalipäivystys (1/1)
uppgjort (1/1)
arbetsintyget (2/2)
studerar (21/21)
då (82/82)
hemförlossning (1/1)
daghemmen (3/3)
vara (146/146)
handlar (2/2)
återflyttning (1/1)
nuorisoasunnot (2/2)
motionsslingorna (1/1)
hindi (1/1)
Itä (1/1)
programmeringsgränssnittfinska (1/1)
utbildats (1/1)
dörrklocka (1/1)
överenskommen (1/1)
Advokatförbunds (1/1)
musik (18/18)
lånet (7/7)
upptäcka (1/1)
brann (1/1)
ögonkontakt (2/2)
universitetens (1/1)
handikappadefinska (3/3)
möjliggör (1/1)
undersökningar (4/4)
underlätta (2/2)
hemkommunens (1/1)
förvärvat (2/2)
beräkning (1/1)
mataffärer (1/1)
begränsa (1/1)
handelstrafik (1/1)
ämnen (10/10)
ärver (2/2)
känslor (1/1)
registret (1/1)
yrkesskolorna (1/1)
swahili (2/2)
bygg- (1/1)
handikappservice (2/2)
valkretsar (1/1)
industriprodukter (1/1)
underhållsstöd (4/4)
flickor (5/5)
grundskolan (33/33)
församlingenfinska (1/1)
förlorar (3/3)
leda (1/1)
vårdar (16/16)
månaderna (5/5)
intagen (1/1)
Ateneum (1/1)
sommarkollon (1/1)
serveras (3/3)
skötaren (2/2)
vigselceremonin (1/1)
delägare (1/1)
Pojkarnas (1/1)
försörja (3/3)
barnatillsyningsmännenfinska (2/2)
biljettjänstens (1/1)
arbetslöshetskassan (6/6)
medlemskortetfinska (1/1)
sambo (17/17)
tjänste- (1/1)
kraftiga (1/1)
förlossningsdatumet (3/3)
natten (2/2)
fritid (4/5) Fritid (1)
skolpsykologen (2/2)
aluekoordinaattori (2/2)
poliisi (1/1)
kraft (13/13)
besiktningskontor (1/1)
samborna (3/3)
kväv (1/1)
konsertsalar (1/1)
Brottsofferjourens (2/2)
pojkens (1/1)
rekryteringen (1/1)
billigare (2/2)
vårdkostnadsförsäkring (1/1)
Uskonnot (2/2)
biljetten (1/1)
behovet (6/6)
preventivmedelsrådgivningens (1/1)
eftersom (19/19)
metron (2/2)
ammatillinen (3/3)
än (106/106)
kinesiska (36/36)
färdigheter (22/22)
ändras (4/4)
psykoterapifinska (1/1)
tidsbundet (7/7)
hälsocentralen (2/2)
naturskyddsområde (2/2)
sidan (36/36)
överbefälhavare (1/1)
storprojekt (1/1)
invandrarkvinnor (10/10)
givet (1/1)
festivaler (1/1)
makan (8/8)
mentalvårdstjänsternafinska (1/1)
sätter (2/2)
grund- (1/1)
anvisningar (19/19)
flyktingläger (2/2)
adresser (3/3)
gäst (2/2)
runtom (3/3)
www.infofinland.fi (1/1)
ansökningsbilagorna (6/6)
färdas (4/4)
VR (1/1)
verkställande (1/1)
nivåerna (2/2)
mobbad (1/1)
hälsovårdsstationen (1/1)
jordbruk (1/1)
intressen (7/7)
kanaler (5/5)
gymnasiekurser (1/1)
ammattitutkinto (1/1)
orättvist (1/1)
utvecklingsstörningar (1/1)
slott (4/4)
utbud (1/1)
flyttsak (2/2)
lekens (1/1)
ansökningsprocessen (1/1)
skäliga (4/4)
EMMAfinska (1/1)
godkänt (4/4)
automatiskt (7/7)
innerstad (1/1)
telefonabonnemang (1/1)
hyresvärd (2/2)
försäljningsmetoder (1/1)
tror (2/2)
flesta (29/29)
kultur (13/13)
ting (3/3)
ord (4/4)
högutbildade (1/1)
LinkedIn (1/1)
kristelefonfinska (1/1)
asylsökande (22/22)
modern (20/20)
isdubbar (1/1)
isär (3/3)
vak (1/1)
bytas (1/1)
spårvagnar (1/1)
frispråkighet (1/1)
parkeringsavgiften (1/1)
uppehållskortet (3/3)
bemötts (1/1)
ena (16/16)
Kelviå (5/5)
arbetarskyddsmyndigheter (1/1)
oikeus (1/1)
specialfall (1/1)
tillbringa (1/1)
grundundervisningenfinska (1/1)
ekonomiplaneringen (1/1)
lagt (1/1)
integrationsåtgärderna (1/1)
yhdistys (1/1)
skolåldern (21/21)
uppväxtmiljö (1/1)
uppenbart (1/1)
stiftelser (3/3)
yläkoulu (1/1)
hotat (2/2)
Korkalovaara (1/1)
ingen (22/22)
sexåringar (2/2)
ungerska (8/8)
kristendomen (1/1)
översättningstjänsterfinska (1/1)
Schengenområdet (6/6)
klubbar (6/6)
barnen (25/25)
övervaka (1/1)
invandrarbyrå (2/2)
kranvatten (1/1)
mitten (3/3)
hinder (15/15)
arbetslösa (25/25)
välja (16/16)
toleransen (1/1)
kaupunginvaltuusto (1/1)
olaglig (1/1)
Runeberg (1/1)
slutar (9/9)
Yhden (2/2)
utbildnings- (1/1)
moder (1/1)
förråd (1/1)
internationell (2/3) Internationell (1)
kapital (2/2)
kunskaper (27/27)
landskapsplanerare (1/1)
konst- (1/1)
flest (2/2)
stödcentret (3/3)
högskolestuderandefinska (1/1)
surfplattan (1/1)
assistans (1/1)
aikuislukio (4/4)
ungdomarnas (2/2)
textning (1/1)
befrämjande (1/1)
uppges (3/3)
sjuksköterska (2/2)
specialbibliotek (1/1)
behandlats (1/1)
vattenånga (1/1)
uppmärksammar (1/1)
vikens (1/1)
demokrati (1/1)
arbetskamraterna (1/1)
sjukvårdsersättningar (1/1)
serviceställena (1/1)
sairaalan (1/1)
besvärlig (1/1)
vammaistuki (2/2)
lilla (1/1)
självständigheten (1/1)
Fernissan (1/1)
industrialisering (1/1)
världen (2/2)
påsk (1/1)
fakulteten (1/1)
handling (4/4)
kliniker (2/2)
företagsverksamhet (15/15)
lånekort (1/1)
lånekostnaderna (1/1)
umgängetfinska (1/1)
mindre (24/24)
ta (117/117)
samlas (3/3)
skatten (2/2)
medarbetare (1/1)
funktionell (1/1)
Barnkliniken (3/3)
gränssnittetfinska (1/1)
eventuellt (11/11)
anställningsrådgivningen (1/1)
gemensamma (37/37)
tusentals (2/2)
handikapprådgivningen (2/2)
aktier (2/2)
försäkringsbolag (11/11)
skriva (16/16)
spelproblemfinska (1/1)
studiemetoder (1/1)
jobbsökning (4/4)
intelligenta (1/1)
tjänstekollektivavtal (1/1)
giftorätt (1/1)
tolkningen (8/8)
helgdag (1/1)
startande (1/1)
stödpersoner (1/1)
bruksföremål (1/1)
A2.1 (1/1)
kartong (1/1)
fullgjorts (2/2)
present (1/1)
egendomen (16/16)
par- (1/1)
sommaruniversitetets (1/1)
ungdomen (1/1)
viss (20/20)
ordningsnumret (1/1)
kunnallisvaalit (1/1)
kontaktperson (1/1)
krissituationer (8/8)
bedömer (16/16)
Omnia (3/3)
försvunnit (1/1)
skickas (8/8)
Silkesportens (1/1)
Indien (1/1)
mobil (1/1)
okomplicerat (1/1)
minska (1/1)
trafikförbindelser (1/1)
bra (54/54)
säsongsarbetefinska (1/1)
sorteras (1/1)
förlossningsavdelningen (1/1)
fri (1/1)
hyra (21/21)
sammankallas (1/1)
gruppfamiljedaghem (4/4)
delta (35/35)
presidentval (4/4)
maximitiden (1/1)
rusmedelsbruk (1/1)
leva (6/6)
intressebevakningsorganisationer (1/1)
rundvandringar (2/2)
aktiivimalli (1/1)
bilaga (1/1)
besluten (1/1)
språkexamen (10/10)
symptom (2/2)
biografen (1/1)
såväl (5/5)
-lokaler (1/1)
speciell (2/2)
stärka (1/1)
skrivit (1/1)
stilla (1/1)
vanligaste (8/8)
bolagsmannen (1/1)
begravningsplats (8/8)
besökarna (1/1)
examensdel (2/2)
datum (2/2)
försäljningen (4/4)
hälsovårdsverket (1/1)
hyresförhållandet (2/2)
A2 (2/2)
självständighet (2/2)
stadsrättigheter (1/1)
måndagar (3/3)
faderskapet (12/12)
socialarbetare (10/10)
genomgår (1/1)
Ab (2/2)
läkemedlen (1/1)
identitetskort (7/7)
städer (22/26) Städer (4)
pappret (1/1)
Pääkaupungin (2/2)
omständighet (1/1)
spisfläkten (1/1)
säsongsarbetstillstånd (1/1)
livscykel (1/1)
läsesal (1/1)
transformera (1/1)
linkkiMiljöministeriet (1/1)
kopiera (2/2)
kallad (2/2)
skrift (1/1)
seger (1/1)
skolbarnfinska (3/3)
plastförpackningar (1/1)
återkalla (1/1)
G (1/1)
anställningar (4/4)
hävas (2/2)
biblioteket (17/17)
pappaledig (1/1)
bekostar (1/1)
lottar (1/1)
arbetskraftsutbildningfinska (1/1)
utser (3/3)
läkaren (20/20)
medicineringen (1/1)
våning (4/4)
befann (1/1)
reklammedel (1/1)
församlingarfinska (1/1)
Linja (7/10) linja (3)
strejk (1/1)
numret (9/9)
arbetar- (1/1)
vårdnadshavare (23/23)
språkkursernas (1/1)
utbildningens (1/1)
stödfunktioner (1/1)
förmånligare (9/9)
begåtts (2/2)
bekant (2/2)
innehar (2/2)
erövrats (1/1)
adoption (3/3)
utlåtande (9/9)
litar (1/1)
former (4/4)
bodelningsman (2/2)
samtalshjälp (4/4)
branschspecifika (1/1)
världsarven (1/1)
arbetsgivares (1/1)
laitos (2/2)
utkomststödfinska (1/1)
anslutna (1/1)
legalisering (2/2)
språk (85/85)
upplösande (1/1)
servicepunkt (1/1)
rättsliga (1/1)
mottagning (4/4)
sönder (1/1)
förstörs (2/2)
kt (5/5)
sträcker (1/1)
frihet (1/1)
Kunta (5/5)
kristen (1/1)
anställningsavtalets (1/1)
Nuppi (3/3)
utkomstskydd (9/11) Utkomstskydd (2)
arbetslöshetsstöd (1/1)
Metropolia (1/1)
flyktingarfinska (3/3)
län (3/3)
fritt (14/14)
senare (11/11)
tandklinik (4/4)
populära (4/4)
integrationsplanfinska (1/1)
situationerna (1/1)
studiemiljön (1/1)
delägarbostadfinska (2/2)
människohandel (12/12)
torka (1/1)
pappersrecept (1/1)
universitetetfinska (1/1)
utövar (7/7)
språkkunskapskrav (1/1)
2:a (1/1)
seniorerfinska (1/1)
turistbyrån (1/1)
makarfinska (1/1)
telefonledes (4/4)
arbets- (58/59) Arbets- (1)
döms (1/1)
skadegörelse (1/1)
hemsidor (2/2)
utbildar (2/2)
peruskielitaito (1/1)
motionsplatserna (1/1)
beträffande (2/2)
styrelse (2/2)
sopbehållare (1/1)
symtomen (1/1)
Virtanen (2/2)
ärva (2/2)
förhistoria (1/1)
överlåtelseskatt (3/3)
samtalsstöd (1/1)
fordonfinska (1/1)
driftställe (1/1)
igenom (5/5)
universitetscenter (1/1)
inkorporerades (1/1)
huvudsyssla (3/3)
pääkaupunkiseudun (1/1)
sysselsättningsplan (4/4)
yrke (16/16)
käpp (1/1)
latauspiste (1/1)
matfinska (1/1)
Vasagatan (1/1)
vigseln (9/9)
utnyttja (13/13)
likaberättigandefinska (1/1)
leder (8/8)
mångsidigt (1/1)
opiskeluterveydenhoitajat (1/1)
Optia (1/1)
nya (40/40)
arbetsför (1/1)
hjälpmedlen (2/2)
domstolsbeslut (4/4)
hyresbostäderfinska (5/5)
sällskapande (3/3)
tiderna (1/1)
att (1223/1233) Att (10)
diskutera (7/7)
tors (5/5)
tjänstens (2/2)
pauser (2/2)
finlandssvenska (2/2)
upprättat (3/3)
kostnader (9/9)
smittsamma (2/2)
kvällstid (4/4)
underleveransarbete (1/1)
Museiverkets (2/2)
natt (1/1)
jourmottagningen (17/17)
därifrån (1/1)
farfinska (1/1)
förhandsröstningsställe (1/1)
umgås (1/1)
tidsbeställningen (2/2)
obegränsad (2/2)
oppisopimus (1/1)
försiktig (1/1)
Novgorod (2/2)
tullanmälan (1/1)
elvärme (1/1)
glasögon (1/1)
förvaltningen (2/2)
skadats (4/4)
filmvisningar (1/1)
skyddar (1/1)
kurserna (16/16)
barnet (160/160)
samorganisation (1/1)
familjens (21/21)
Myrbackahuset (1/1)
kursstart (1/1)
psykoterapeutti (1/1)
flytväst (1/1)
familjebostäder (1/1)
vet (6/6)
Saarnio (2/3) saarnio (1)
sjukt (6/6)
stärker (1/1)
hemsida (1/1)
indoeuropeiska (1/1)
myndighet (11/11)
rekreation (1/1)
augusti (6/6)
inträdesprovet (2/2)
flygeln (1/1)
deltid (5/5)
reserverad (1/1)
könsidentitet (3/3)
yrkeshögskolekurser (1/1)
placeras (1/1)
Vantaan (10/10)
framtidens (1/1)
folkhögskola (2/2)
arabiska (59/59)
recept (15/15)
tandvården (6/6)
respekteras (1/1)
långvarigt (1/1)
studieområde (1/1)
asuminen.fifinska (2/2)
RAOS (1/1)
nödnumret (32/32)
garantipensionerna (1/1)
borgensmän (1/1)
ambulans (1/1)
arbetsolycksfall (1/1)
kommanditbolaget (1/1)
uppehållstillståndsärenden (1/1)
läroavtalscenterfinska (1/1)
Omatila (4/4)
integritet (3/3)
innehållits (1/1)
nybörjareengelska (1/1)
befogade (1/1)
finansiering (12/12)
bekantat (1/1)
när (196/202) När (6)
avgörs (1/1)
upphörde (1/1)
sö (1/1)
Health (1/1)
droger (5/5)
journumret (2/2)
plastföremål (1/1)
ryssarna (1/1)
egnahemshuset (1/1)
Nuortennettifinska (1/1)
räknats (1/1)
förlikning (2/2)
stadsbibliotek (7/7)
tio (3/3)
meddelanden (1/1)
inlärningsgrupp (1/1)
minnestest (1/1)
konsumenträttigheterfinska (1/1)
har (1057/1057)
makes (5/5)
barnklubbar (3/3)
servicestället (10/10)
bortfaller (1/1)
talets (1/1)
förts (1/1)
tjeckiska (1/1)
ställena (1/1)
uppehälle (5/5)
babyn (3/3)
integration (13/18) Integration (5)
ovanför (2/2)
främjande (2/2)
chefer (1/1)
hans (10/10)
kielitaito (2/2)
barnatillsynsmannen (1/1)
K.H.Renlunds (3/3)
skriver (11/11)
bankärendenfinska (1/1)
glaset (1/1)
grannmedlingscentret (1/1)
täcker (3/3)
lägre (9/9)
april (4/4)
tidsbeställning (7/7)
sommaruniversitetfinska (2/2)
någonstans (3/3)
gammal (13/13)
Axxell (2/2)
stiftelsen (2/2)
exceptionellt (2/2)
harkinnanvarainen (1/1)
musikundervisning (1/1)
brandlarm (1/1)
gymnasieböckerna (3/3)
uppehållskort (5/5)
hus (7/7)
aborten (1/1)
uppehållstillståndet (14/14)
högskolor (12/13) Högskolor (1)
ägande (1/1)
invånarantalet (1/1)
turistersvenska (1/1)
likadant (1/1)
behandlingsmetoder (1/1)
morbror (1/1)
AUS (1/1)
registrerats (3/3)
hålla (4/4)
hyreslägenheten (1/1)
integrationsutbildningen (2/2)
C1 (1/1)
Verso (1/1)
skolans (10/10)
sexuellt (7/7)
mångfaldigades (1/1)
bebiskläder (1/1)
bedöma (3/3)
ungdomsbostäder (5/5)
innanför (1/1)
lampa (1/1)
kroppsaga (2/2)
välityspalkkio (1/1)
innehåll (5/5)
redaktion (2/2)
avstå (1/1)
kursen (4/4)
stadsfullmäktige (7/7)
åtalas (1/1)
faderskapsledigheten (3/3)
gym (3/3)
högskoleexamen (18/18)
grannen (1/1)
problematiskt (1/1)
församlingfinska (1/1)
myndighetstjänst (1/1)
invandrarmän (3/3)
diskriminering (37/39) Diskriminering (2)
vigseltiden (1/1)
anställningsavtal (1/1)
utöver (5/5)
Kristinestad (1/1)
montera (1/1)
settlementföreningen (1/1)
rabatter (1/1)
byggherrar (1/1)
hyresgarantin (2/2)
accepterade (1/1)
asylsamtal (1/1)
rad (1/1)
luftfartsyrken (1/1)
Muurola (1/1)
bokhandlar (1/1)
hyresboendefinska (1/1)
specifikationsdel (2/2)
partnerskap (2/2)
positivt (4/4)
läroavtalscenter (3/3)
egendom (28/28)
huvudsakliga (1/1)
underlättar (6/6)
justitieministeriets (2/2)
etablerades (2/2)
fågelbon (2/2)
tolkcentral (3/3)
finnas (10/10)
begravningfinska (1/1)
kopplas (2/2)
dagtid (3/3)
förgiftningfinska (1/1)
Elfvik (1/1)
affärspartner (1/1)
förnya (4/4)
Clinicin (1/1)
hushållsmaskin (1/1)
under (232/232)
bassjälvrisken (1/1)
Espoon (7/7)
flyttar (86/86)
juni (9/9)
återkallats (2/2)
överlåtelse (1/1)
snabbköp (1/1)
användas (6/6)
hälsotjänsterna (3/4) Hälsotjänsterna (1)
yttranderätt (1/1)
kontrolleras (3/3)
någons (1/1)
föreskrivas (1/1)
redovisning (2/2)
linje (2/2)
hushållsapparater (1/1)
oavbrutet (1/1)
Sanduddsgatan (1/1)
grundtryggheten (1/1)
kriisipalvelu (1/1)
verifieras (1/1)
gonorré (1/1)
vuxenutbildningsstöd (1/1)
prövning (11/13) Prövning (2)
övertidsarbete (1/1)
pojkvän (1/1)
erbjuder (79/79)
Kylämajafinska (1/1)
nätbankskoderna (1/1)
tilläggsstudier (1/1)
vatten (4/4)
församlingssammanslutnings (2/2)
anordnad (2/2)
vårdledig (3/3)
germanska (1/1)
työttömyyskassa (1/1)
linjen (1/1)
seniorrådgivning (1/1)
farligt (4/4)
startpenning (5/5)
byråfinska (1/1)
skattemedel (1/1)
region (2/2)
guidar (1/1)
ger (82/83) GER (1)
kvarskatten (1/1)
organen (1/1)
begravningsbyråer (2/2)
kirkko (2/2)
utöka (2/2)
familjeträningen (1/1)
familjebandfinska (2/2)
du (2752/2757) Du (5)
Nuorisoasiainkeskus (1/1)
ändamål (1/1)
Kiinteistöyhtiö (1/1)
Finnish (2/2)
fyller (17/17)
företagarefinska (6/6)
klinikens (5/5)
högskolornas (3/3)
döva (1/1)
skör (1/1)
myndiga (2/2)
invånarinitiativ (1/1)
ert (1/1)
jobbsökningenfinska (1/1)
fysiskt (1/1)
Navigatorn (5/5)
ledamöterna (1/1)
lapsilisä (1/1)
Apotekareförbundets (1/1)
program (8/8)
lämna (39/39)
österifrån (1/1)
begravas (3/3)
identitetsnummer (1/1)
behandlingen (7/7)
livssituation (7/7)
medborgarnas (2/2)
ansöks (4/4)
räcker (11/11)
hoidon (1/1)
palvelu (1/1)
oumbärliga (1/1)
tåg (3/3)
upphör (18/18)
empirestil (1/1)
tjänstebehörighet (2/2)
skolor (18/18)
hyreskontrakt (2/2)
relaterade (1/1)
nej (1/1)
kristna (3/3)
styrs (2/2)
biograf (2/2)
äktenskapfinska (2/2)
språkkunskapskraven (1/1)
sjukförsäkring (8/8)
arbetsintygfinska (1/1)
maksuhäiriömerkintä (1/1)
viitekehys (1/1)
telefonabonnemangfinska (1/1)
kallelse (1/1)
hota (1/1)
klienten (2/2)
framgå (3/3)
bedrevs (1/1)
skilsmässoansökan (6/6)
likvidation (1/1)
medlemmarna (3/3)
makens (4/5) Makens (1)
intressant (2/2)
anvisa (1/1)
tillgodoräknas (2/2)
antecknas (4/4)
förfallodagen (2/2)
examenstillfällen (1/1)
sökas (4/4)
finnishcourses.fi (2/4) Finnishcourses.fi (2)
vidimera (1/1)
underhållsskyldighet (2/2)
välbefinnandet (1/1)
antas (3/3)
vederbörliga (2/2)
julen (2/2)
servicenivån (1/1)
föreläsningsserier (1/1)
farföräldrarna (1/1)
registrering (20/29) Registrering (9)
betyg (4/4)
buffert (1/1)
integrationsplan (14/14)
videoklipp (3/3)
Vanhemman (2/2)
barnlösheten (1/1)
kartanfinska (1/1)
pensionering (1/1)
arbetarskyddsdistriktet (1/1)
Sinettä (1/1)
vårdanstalter (1/1)
förhandla (2/2)
lukiopohjainen (1/1)
visst (6/6)
förbereds (1/1)
faderns (4/4)
beroendeproblem (1/1)
gårdsområden (1/1)
Eija (2/2)
kista (1/1)
använd (2/2)
framhävs (2/2)
studiestödetfinska (1/1)
skatteprocenten (2/2)
betjänas (1/1)
Vanttauskoski (1/1)
alkoholisterfinska (1/1)
hanke (1/1)
konventionsstaterna (1/1)
åring (1/1)
säsongtopp (1/1)
areal (3/3)
hand (60/60)
levereras (1/1)
vända (7/7)
människa (2/2)
livmoderns (1/1)
Punaisen (2/2)
idrottsområdet (4/4)
privatsfär (1/1)
finskakurser (3/3)
Konvaljvägen (1/1)
Isyysraha (1/1)
työsuojelupiiri (1/1)
Anders (1/1)
röstning (2/2)
främst (5/5)
missbrukarefinska (2/2)
arbetslöshetsförmånerfinska (1/1)
uppsöka (1/1)
språktest (1/1)
vårdpenning (10/10)
företagsform (2/2)
kyrkan (21/21)
E101 (2/2)
Noux (1/1)
smidigt (1/1)
krismottagning (2/2)
invandrarbyrån (4/4)
lämplig (14/14)
kallade (3/3)
genomtänkta (1/1)
förhållanden (2/2)
bolagsvederlag (1/1)
resmålet (1/1)
åker (5/5)
regionutvecklingen (1/1)
filosofi (1/1)
trupper (1/1)
festlokal (1/1)
bostadsvisning (2/2)
patientavgift (1/1)
roliga (1/1)
ansikte (2/2)
kyrka (5/5)
rekommendera (2/2)
skatteförvaltningenfinska (1/1)
instans (3/3)
Olkkarifinska (1/1)
-eller (1/1)
doulaverksamheten (1/1)
myhelsinki.fi (1/1)
oavsett (7/7)
underhåll (5/5)
hamnade (1/1)
info (8/8)
räknas (10/10)
biograferna (1/1)
uppdatera (2/2)
individualism (1/1)
finländsk (18/18)
faderskapsärendet (1/1)
parter (1/1)
nackdel (1/1)
klarläggs (1/1)
kravet (3/3)
sökfunktionen (1/1)
helsingforsare (1/1)
Vandas (2/2)
rekommendationer (1/1)
utbildning (87/92) Utbildning (5)
kassan (5/5)
snittbetyg (1/1)
avgångsbetyg (5/5)
servicenumret (1/1)
skadas (1/1)
teckenspråket (1/1)
Vionojas (1/1)
oss (1/1)
tilläggsdagar (1/1)
beskattningsbeslut (1/1)
skogsbruksingenjör (1/1)
hamnverksamheten (1/1)
lasi (1/1)
låneräknare (1/1)
stängt (6/6)
miljöer (1/1)
tidningarna (1/1)
responslänk (1/1)
FPA (94/108) Fpa (14)
språkkaféerna (1/1)
låga (4/4)
työväenopisto (4/4)
socialarbetaren (2/2)
individuellt (3/3)
boendefinska (1/1)
hälsovårdsenhet (1/1)
påverka (25/25)
skilsmässan (5/5)
studerande (52/54) Studerande (2)
intressebevakningsorganisationfinska (1/1)
inlärningen (1/1)
bild (2/2)
ständigt (1/1)
länder (36/36)
handarbeten (3/3)
giltig (2/2)
läroanstalterna (2/2)
kroatiska (4/4)
inredningsarkitekt (1/1)
sommargymnasium (1/1)
fågelungar (2/2)
barnskyddslagen (1/1)
förplikta (1/1)
besöksförbudfinska (1/1)
förorter (1/1)
centralernafinska (1/1)
typen (1/1)
rådgivningsbyråerna (3/3)
växer (2/2)
varierande (1/1)
avbokat (1/1)
brott (48/50) Brott (2)
Estnäs (1/1)
åtgärder (4/4)
vartannat (3/3)
urologiska (1/1)
klara (16/16)
handikappidrott (1/1)
både (24/24)
rättshjälpsbyråer (1/1)
elbolag (1/1)
rehabiliteringsplan (2/2)
förmyndarskap (2/2)
måla (1/1)
tryggar (8/8)
flyktingstatus (16/16)
elever (9/9)
integrationsstöd (1/1)
tycker (1/1)
vårdnadshavarna (2/2)
skyldigheterfinska (1/1)
Utbildningsstyrelsens (13/17) utbildningsstyrelsens (4)
parken (1/1)
vårdnadshavaren (1/1)
urvalsbaserade (1/1)
avgöras (1/1)
tjänsteman (1/1)
ofött (1/1)
heltidsstudier (4/4)
Nordplus (1/1)
tillsammans (56/56)
Jesu (3/3)
Giftinformationscentralen (1/1)
antecknar (1/1)
regionkontorfinska (1/1)
kraven (2/2)
förknippade (2/2)
kopior (2/2)
vintrarna (1/1)
plötsliga (1/1)
industrialiseringen (2/2)
startpengen (1/1)
vuxengymnasierna (1/1)
sön (2/2)
roligt (1/1)
uppgifterfinska (1/1)
Oulun (1/1)
resorna (1/1)
Laurea (2/2)
förutsatt (1/1)
café (1/1)
postfinska (1/1)
torteras (1/1)
bibliotekarienfinska (1/1)
Alkoholistit (1/1)
dra (3/3)
arbetskraft (2/2)
päivystysajanvaraus (1/1)
högstadiet (4/4)
beslutsfattande (3/3)
byrån (54/54)
hennes (9/9)
valdagen (8/8)
övergår (1/1)
pågår (16/16)
stödboende (3/3)
debiteras (1/1)
registrerades (2/2)
läroanstalten (11/11)
översättar- (3/3)
rättshjälpfinska (1/1)
nationellt (1/1)
andel (6/6)
uträttar (3/3)
privat (46/46)
eläkekassa (1/1)
orten (4/4)
handelsflotta (1/1)
begår (4/4)
Sello (1/1)
familjer (25/28) Familjer (3)
mödrahemmet (2/2)
avslag (2/2)
bastuugnen (3/3)
parkerna (1/1)
Al (1/1)
ammattikorkeakoulututkinto (1/1)
öppettiderfinska (2/2)
kerho (1/1)
förskoleundervisningen (13/13)
sosiaaliohjaaja (1/1)
Religionerna (1/1)
undervisningsväsendet (1/1)
lagar (13/13)
invandrarföreningar (3/3)
ombud (1/1)
arbetskraftsutbildningen (2/2)
kommunikationssvårigheter (1/1)
breddgraderna (1/1)
Karlebys (2/2)
sorg (1/1)
doktorsexamen (4/4)
begravningsplatsfinska (1/1)
yrket (1/1)
vetenskapsbibliotek (1/1)
lantdag (1/1)
når (1/1)
butiker (2/2)
modersmålsprovet (2/2)
rättvist (3/3)
Kalkkers (1/1)
invandrarbarn (4/4)
hälsovårdare (19/19)
kulturcentral (1/1)
Utbildningsstyrelsen (3/3)
begagnade (1/1)
olycka (10/10)
verksamhetsspråk (1/1)
hör (26/26)
bestämmer (4/4)
rekisterihallitus (1/1)
förmögenhet (3/3)
århundradet (1/1)
etc (1/1)
förbindelse (2/2)
hemlandet (2/2)
arbetskraftsmyndigheten (1/1)
kielitutkinto (3/3)
yliopistollinen (1/1)
miljön (3/3)
fördröjas (1/1)
överväger (7/7)
socialjouren (2/2)
återvändande (1/1)
reglerar (1/1)
bouppteckningfinska (1/1)
bedömningar (1/1)
hyresbeloppet (1/1)
vetenskaps- (3/3)
bilens (1/1)
Oma (1/1)
varandra (16/16)
beskrivs (2/2)
Galoppbrinken (1/1)
sommaruniversitet (2/2)
godkännande (1/1)
fungerande (1/1)
avgiftsfri (10/10)
listan (2/2)
licentiat- (1/1)
nämnden (1/1)
tjänat (1/1)
förvärvsarbete (2/2)
ambassad (1/1)
alkukartoitus (2/2)
gravida (8/8)
bostadsrättsavgiften (4/4)
böjs (2/2)
lag (37/37)
centrum (9/9)
hanteras (2/2)
personerfinska (1/1)
dörrar (1/1)
betänketiden (5/5)
ring (10/12) Ring (2)
fackförbundet (5/5)
Vuxeninstitut (1/1)
besiktningsstationer (2/2)
folkpensionerna (1/1)
födseln (4/4)
hälsan (13/13)
ylioppilastutkinto (1/1)
finskakunskaper (1/1)
norra (2/2)
nödsituation (11/11)
boendetid (1/1)
talo (2/2)
läsas (2/2)
framgångsrikt (1/1)
graviditetstest (2/2)
Västra (8/11) västra (3)
tiotusentals (2/2)
tälta (1/1)
dekorerat (1/1)
arbetarskyddsfrågor (1/1)
lediga (12/12)
utbytesprogrammetengelska (1/1)
kansalaisen (1/1)
brottsmålsvittnen (1/1)
bank- (1/1)
Lochteå (1/1)
sjuk (20/20)
existensminimum (2/2)
renoveringen (1/1)
avdrag (5/5)
vakuutus (2/2)
tjänster (128/133) Tjänster (5)
SERI (2/2)
asevelvollisuus (1/1)
vattenkran (1/1)
barnskyddets (2/2)
utrikeshandel (1/1)
normal (2/2)
hämta (6/6)
operationen (5/5)
höstens (1/1)
kommer (62/62)
företagsekonomi (1/1)
studentbostadsstiftelser (1/1)
åldringshem (1/1)
dessa (56/56)
anknytning (2/2)
särställning (1/1)
betalningen (1/1)
kalendermånad (2/2)
ungdomsgrupper (1/1)
nyttig (8/8)
stödhandtag (1/1)
arbetarinstitutens (1/1)
tillträde (2/2)
responsiv (1/1)
Kampen (2/2)
evankelis (1/1)
matkakortin (1/1)
angående (3/3)
nödvändigtvis (10/10)
hälsa (63/69) Hälsa (6)
trygghetfinska (1/1)
skador (3/3)
handelsregistret (2/2)
sökanden (3/3)
avgift (2/2)
cykel- (1/1)
kesäyliopisto (1/1)
lönetillägg (1/1)
hemvårdsstödets (1/1)
apparater (2/2)
sjunde (1/1)
jourtelefon (1/1)
ibruktagande (1/1)
stöd- (2/3) Stöd- (1)
undgår (1/1)
himmelsfärd (1/1)
revisionsbyrå (1/1)
uppehållsrätt (28/28)
To (4/4)
lista (7/9) Lista (2)
samlats (1/1)
ryskspråkiga (1/1)
kommunikationen (1/1)
lämnat (3/3)
förmånen (1/1)
uppehållstillståndetfinska (1/1)
voimavarakeskus (1/1)
tidningsannonser (2/2)
blivande (3/3)
dagliga (12/12)
arbetstiden (4/4)
Commons (1/1)
folkpensionen (1/1)
nattjour (3/3)
spel (4/4)
lån (23/23)
avlägger (10/10)
miljö (5/5)
störa (1/1)
matkulturer (1/1)
ledig (1/1)
teckna (9/9)
lagman (1/1)
anger (3/3)
ovanligt (1/1)
sederengelska (1/1)
jobb (55/55)
känt (1/1)
Pakolaisneuvonta (2/2)
följs (11/11)
föräldraledig (3/3)
stadissa.fi (2/2)
invånarna (10/10)
Baltikum (1/1)
fåglar (1/1)
studiepenningen (1/1)
drogmissbruk (1/1)
familjeverksamhet (1/1)
sinsemellan (1/1)
helsinki.fi (1/1)
andelslaget (1/1)
finskspråkiga (14/14)
barnmorska (1/1)
efternamnet (2/2)
diskrimineringsfall (1/1)
experterna (1/1)
äts (1/1)
bostadsrättsbostad (10/11) Bostadsrättsbostad (1)
mossa (1/1)
arbetarskyddsfullmäktige (2/2)
förlängd (1/1)
kaikille (1/1)
tilläggsinformation (1/1)
etälukio (1/1)
slags (17/17)
kypsyysnäyte (1/1)
företett (1/1)
diskrimineringsombudsmannen (2/3) Diskrimineringsombudsmannen (1)
familjepensionfinska (1/1)
hemvårdsstödfinska (2/2)
uppgå (2/2)
närbibliotek (1/1)
avlider (4/4)
längden (1/1)
medlemskap (2/2)
helgdagar (4/4)
antecknats (3/3)
hemspråksundervisningfinska (1/1)
24h (3/3)
rättsbiträde (3/3)
statsöverhuvud (1/1)
intygen (1/1)
synskadade (4/4)
själva (12/12)
misstänker (11/11)
läkarundersökning (4/4)
funderar (5/5)
förtjänat (1/1)
läkemedel (25/29) Läkemedel (4)
skilt (3/3)
fenomen (1/1)
hemkommunfinska (1/1)
ryska (146/146)
invalidpension (4/4)
mental (8/9) Mental (1)
kontor (4/4)
håll (10/10)
partier (1/1)
teater (8/8)
navigator (1/1)
Enter (26/26)
FRK (1/1)
förs (3/3)
mentor (2/2)
tillslutas (1/1)
freelancer (1/1)
invandrarkvinnorfinska (1/1)
Fulbright (2/2)
arbetsdagen (2/2)
-stiftelser (1/1)
svag (1/1)
ämbetsverk (1/1)
tecknar (2/2)
genomförs (2/2)
unionens (2/2)
Europafinska (1/1)
hotell (1/1)
västerut (1/1)
allaktivitetscentret (1/1)
invandrarefinska (20/20)
fängelsestraff (3/3)
kortfinska (1/1)
Nylandfinska (1/1)
inledningsvis (1/1)
BY (2/2)
säkerhets- (1/1)
forststyrelsens (1/1)
Terveyden (1/1)
servicebostäder (1/1)
hallitus (1/1)
lääkinnällinen (1/1)
barnfamiljerfinska (2/2)
studiekamrater (1/1)
månader (71/71)
tiotals (1/1)
royaltyn (1/1)
ungdomslokalerna (1/1)
koulumatkatuki (1/1)
bolagets (1/1)
försöker (6/6)
bostad (102/102)
industri (2/2)
centrala (8/8)
flygplatser (1/1)
House (2/2)
skuldrådgivare (1/1)
ersättning (16/16)
företagande (12/12)
grunden (5/5)
begravningsbidrag (1/1)
riksdagens (1/1)
svenskspråkig (8/8)
åkrarna (1/1)
hälso- (20/20)
utbetalning (4/4)
skattebyrån (13/13)
världsarv (2/2)
bostadslånfinska (1/1)
uppgiften (3/3)
själv (93/93)
felaktiga (3/3)
pensionstagarefinska (1/1)
mångfacetterad (1/1)
skattepliktiga (1/1)
välmående (3/3)
regeringarna (1/1)
varieteter (1/1)
årfinska (2/2)
familjerådgivningscentral (3/4) Familjerådgivningscentral (1)
telefonnumren (1/1)
värderingar (1/1)
arbetsförsök (1/1)
älv (1/1)
nordiska (13/13)
kundtjänsten (7/7)
telefonservice (2/2)
tulkkaus (1/1)
handikappservicefinska (4/4)
batterierna (1/1)
yrkeshögskolan (9/10) Yrkeshögskolan (1)
vandra (1/1)
postpositioner (1/1)
källorna (1/1)
A1.3 (1/1)
vardag (2/2)
infektion (1/1)
lokaltrafiken (1/1)
läkarmottagningen (3/3)
missbruksvård (1/1)
arbetslösfinska (1/1)
skyddshemfinska (3/3)
ersatts (1/1)
älvar (1/1)
inom (99/99)
arbetsplatsens (4/4)
kvinnor (34/34)
uppträder (2/2)
förövaren (1/1)
skogsmuseumfinska (1/1)
lämplighetsprov (1/1)
beslutet (13/13)
avbryts (3/3)
husdjur (1/1)
albanska (7/7)
Startup (1/1)
börjat (3/3)
penningbelopp (1/1)
redaktionen (1/1)
köpebrevet (1/1)
illegala (1/1)
storstäderna (1/1)
vändagen (2/2)
rådgivningsbyråer (6/6)
insjukna (1/1)
utexamineras (1/1)
vanlig (3/3)
etableringsanmälan (2/2)
familjerådgivningscentralen (1/1)
ansökanfinska (2/2)
delägarbostäder (4/4)
giltighetstiden (2/2)
vindruta (1/1)
handelsmän (1/1)
bostadsaktie (2/2)
läkar- (1/1)
intagna (1/1)
ditt (254/254)
arbetssäkerheten (2/2)
deras (36/36)
följer (12/12)
Uunofinska (1/1)
peruskoulupohjainen (1/1)
omänsklig (1/1)
tillförlitligt (2/2)
kopplat (1/1)
STTK (1/1)
kemikalier (2/2)
lekparkernas (1/1)
slidmynningen (1/1)
bildkonst (8/8)
jobbet (3/3)
besök (8/8)
slutbetyget (1/1)
medborgaren (1/1)
vattenavgift (1/1)
brottsmisstänkta (3/3)
skolkuratorer (1/1)
bostadsbyrå (1/1)
komposteras (1/1)
trygga (8/8)
Dödsfall (1/1)
uppehållstiden (1/1)
hälsorådgivningfinska (2/2)
femton (1/1)
VSB (1/1)
mellanskillnaden (1/1)
specialdagvård (1/1)
marknaden (1/1)
testamentti (2/2)
Tulli (1/1)
nuvarande (7/7)
mognadsprov (2/2)
Ceremonier (1/1)
samarbetsområdet (1/1)
Australien (1/1)
förhand (19/19)
ärenden (58/58)
kulturcentret (1/1)
anställningsvillkoren (2/2)
nationella (2/2)
intagning (1/1)
sparas (2/2)
andelar (1/1)
egenskaperna (1/1)
nedsatt (1/1)
företagskulturen (2/2)
faktiska (1/1)
Olofsborg (1/1)
Karlebystöd (1/1)
försäkringspremier (1/1)
framhäver (1/1)
tredjelandsmedborgare (1/1)
barnpassningshjälpen (1/1)
Yritys (2/2)
skilja (3/3)
specialsmåbarnspedagogiken (1/1)
bokfinska (1/1)
invandrat (2/2)
behärska (1/1)
utgörs (3/3)
kosthållsbranschen (1/1)
dåligt (1/1)
plötsligt (4/4)
Avia (1/1)
sjukledighetsdagen (1/1)
september (3/3)
bli (27/29) Bli (2)
fördelning (2/2)
hälsoundersökning (1/1)
4:e (2/2)
sammanlagt (2/2)
omfattas (43/43)
Ambassader (2/2)
sed (2/2)
pyntas (1/1)
ärlighet (3/3)
cyklister (1/1)
batteri (2/2)
FöPL (1/1)
inhemsk (1/1)
belysta (1/1)
orsaken (6/6)
utträda (1/1)
Naapuruussovittelun (1/1)
invandringsfrågor (1/1)
för- (1/1)
insjuknandet (4/4)
utlänningarfinska (3/3)
utställningarfinska (1/1)
bostadsköpet (1/1)
vuxenutbildningscentra (1/1)
hobbymöjligheterna (1/1)
sent (4/4)
storfurstendöme (1/1)
högskolekoncern (1/1)
WC:n (1/1)
amatörer (1/1)
besöka (35/35)
slå (3/3)
vandring (2/2)
pappa (1/1)
studenthälsovårdarna (1/1)
visum (20/20)
arbetsoförmåga (1/1)
myndigheten (18/18)
beviljas (36/36)
handskar (1/1)
användarpanel (2/2)
dagverksamhet (4/4)
hel.fi (2/2)
förstasida (1/1)
serviceboendefinska (1/1)
avlagda (1/1)
trygg (5/5)
faderlöst (2/2)
oljemängden (1/1)
skyddskårerna (1/1)
kommuns (3/3)
års (16/16)
sevärt (1/1)
Mt (2/2)
krama (1/1)
handlingarna (3/3)
tjänstestället (11/11)
tingsdomare (1/1)
enskilde (1/1)
Kervo (2/2)
beställer (7/7)
klart (1/1)
stadsdirektörer (1/1)
museiområden (1/1)
hemvård (6/6)
förebygga (1/1)
skollov (1/1)
familjedagvården (2/2)
trapphuset (2/2)
rättighet (2/2)
skolbarns (4/4)
djurskötarexamen (1/1)
Kasabergsområdet (1/1)
ateriatuki (1/1)
modersmålsundervisningen (1/1)
ur (8/8)
arrangören (1/1)
gymnasiestudier (6/6)
överens (43/43)
Helsingforsbor (1/1)
obekvämt (1/1)
Fjällrävsstigen (1/1)
perheasioiden (2/2)
föräldraskap (2/2)
sjukförsäkrad (2/2)
biljettpriserna (2/2)
ELY (1/1)
sjukhuset (17/17)
sannolikt (2/2)
hamnar (2/2)
data- (1/1)
besökt (3/3)
Arbetslöshetsförsäkring (5/9) arbetslöshetsförsäkring (4)
rekreationsområde (1/1)
avslår (2/2)
inresereglerna (1/1)
seurakuntien (1/1)
motarbeta (3/3)
Myyrinki (1/1)
tillsyn (1/1)
förhandlar (1/1)
återförening (1/1)
restauranger (1/1)
yleinen (3/3)
armé (1/1)
undersöka (1/1)
tidsbokning (11/11)
Silkinportin (1/1)
motions- (1/1)
elektroniskt (11/11)
samfällighet (3/3)
träffpunkten (1/1)
jämkning (1/1)
seniorrådgivningen (4/5) Seniorrådgivningen (1)
könssjukdomar (8/8)
företagfinska (2/2)
hälsosam (1/1)
mångkulturell (3/3)
vinnare (2/2)
ambassaden (1/1)
fastställande (2/2)
dagligen (1/1)
Mundus (1/1)
företagshälsovården (7/8) Företagshälsovården (1)
yrkesinriktad (31/31)
Ihmiskaupan (1/1)
närståendevåld (1/1)
hyrsvärden (1/1)
undertecknas (1/1)
kotikunta (6/6)
asuntoa (2/2)
slutit (1/1)
stämmor (1/1)
lekparksverksamhetfinska (1/1)
tandläkaren (3/3)
avlidit (1/1)
utvecklades (2/2)
rf:s (3/3)
invånaren (1/1)
börja (16/16)
B1 (2/2)
finländare (11/11)
oftast (22/22)
pengar (10/10)
dåliga (1/1)
linkkiFinnkino (1/1)
förlänga (3/3)
psykoterapin (1/1)
dag (27/27)
firma (1/1)
döda (2/2)
affärsmannen (1/1)
husbolaget (2/2)
hänsyn (5/5)
början (16/16)
gratis (22/22)
tolksbehovet (1/1)
kunder (5/5)
Myrbacka (2/2)
personen (9/9)
sömnskola (1/1)
synagoga (1/1)
tandkirurgi (1/1)
veckoslutet (2/2)
kulturtjänster (2/2)
möblerade (1/1)
registreringsintyg (2/2)
uppriktighet (1/1)
institutets (7/7)
månad (24/24)
loss (1/1)
hyresvärden (18/18)
åringar (5/5)
tryggt (5/5)
åtminstone (13/13)
pojkes (1/1)
regnar (1/1)
handelscentra (1/1)
responssystemfinska (1/1)
farföräldrar (2/2)
böcker (16/16)
vuxensocialarbetetfinska (1/1)
kunnandet (2/2)
nekande (1/1)
erkände (1/1)
diskriminerad (1/1)
utreds (4/4)
återvänder (3/3)
försvunna (1/1)
Tukinainen (1/1)
medverkat (4/4)
muovi (1/1)
ansluter (4/4)
vårt (2/2)
Internetanslutning (1/2) internetanslutning (1)
ansökningstid (1/1)
Arbetseffektivitetsföreningen (2/2)
missgynnas (1/1)
människors (5/5)
arbetarinstitutet (1/1)
Mona (4/4)
läsämnena (1/1)
förvärvsinkomst (2/2)
öppet (38/39) Öppet (1)
lådor (1/1)
ägodelar (2/2)
servicetorget (1/1)
yhdenvertaisuusvaltuutettu (1/1)
uppmuntrar (2/2)
Apteekkariliitto (1/1)
bekräfta (1/1)
skald (1/1)
lyftandet (1/1)
drivas (1/1)
koulunkäyntiavustaja (1/1)
ntresserad (1/1)
bristen (2/2)
skönhetsvård (1/1)
pedagogik (5/5)
oväsen (1/1)
biIdkonstskola (1/1)
vissa (88/88)
relationerna (3/3)
direkt (55/55)
härkomst (4/4)
skiljer (5/5)
guidade (3/3)
familjeskäl (4/4)
Spa (1/1)
ängre (1/1)
testamentsgåva (1/1)
A (25/26) a (1)
mobilcertifikat (3/3)
bestämmanderätt (1/1)
papperspåsar (1/1)
ämnesområden (1/1)
familjeförmånerna (1/1)
avsevärt (3/3)
försvara (2/2)
Vandainfo (1/1)
Asianajajaliitto (1/1)
spelande (3/3)
h (1/1)
Quebec (1/1)
busslinjer (2/2)
familjefrågorfinska (2/2)
avser (6/6)
avtal (30/30)
förtagaren (1/1)
exakt (2/2)
munhälsans (1/1)
videoklippet (12/12)
olika (179/179)
projekt (3/3)
ingås (5/5)
sydkust (1/1)
växa (2/2)
utlandet (13/13)
skoldagen (3/3)
flytta (16/21) Flytta (5)
åren (6/6)
arvo (1/1)
paddlare (1/1)
tågtidtabellerna (1/1)
varat (5/5)
kommit (12/12)
alla (120/120)
huset (4/4)
lunch (3/3)
vecka (7/7)
besöker (10/10)
meritförteckning (5/5)
litet (6/6)
ungdomsstation (1/1)
Poikien (1/1)
medlemsavgift (2/2)
firar (1/1)
utbetalas (9/9)
inslag (1/1)
kostnadsfritt (5/5)
lättföretagande (1/1)
dagar (35/35)
godtar (1/1)
jurist (14/14)
hyresbostadfinska (1/1)
koder (1/1)
Sverige (16/16)
beaktas (14/14)
yrkeshögskolestudier (1/1)
parts (1/1)
krav (4/4)
män (25/25)
uppgett (1/1)
skolresa (1/1)
punkten (1/1)
Arbisfinska (1/1)
förmedlingsarvodet (3/3)
mössa (1/1)
närmast (5/5)
helhetsbetonat (1/1)
kierrätyspiste (1/1)
visumcentral (1/1)
arbetsplatser (13/13)
barnfostran (1/1)
studentexamen (7/7)
inskolning (3/3)
väntar (6/6)
avtala (1/1)
framgår (3/3)
pappersblanketter (1/1)
hälsorådgivningens (1/1)
tingsrätts (2/2)
poliklinikka (3/3)
anvisar (2/2)
beskriver (5/5)
caféerna (1/1)
veckan (4/4)
försvarandet (1/1)
Caisa (1/1)
Sporttia (1/1)
utfärda (6/6)
avslutas (1/1)
exakta (3/3)
förbundets (2/2)
bestraffas (1/1)
skenäktenskap (1/1)
diskussioner (2/2)
konfessionslösa (2/2)
tuki (5/5)
tillhandahålla (2/2)
skrapning (2/2)
Domus (1/1)
flytt (8/8)
arbetssäkerhets- (1/1)
Kehitysvammahuollon (1/1)
byarna (1/1)
må (1/1)
språkexaminafinska (4/4)
motionsdosen (1/1)
kyrkliga (5/5)
bastuugn (2/2)
färdig (1/1)
tidtabellerfinska (1/1)
Rovalas (1/1)
giftorätten (1/1)
turvakaukalo (1/1)
vårdare (1/1)
Väestöliitto (6/6)
sammanslutning (1/1)
höja (4/4)
nyföretagarcentralerna (1/1)
integrationsplanen (9/9)
studiekraven (1/1)
samhällsgrupp (2/2)
psykiater (1/1)
råder (2/2)
mathjälp (1/1)
högskolan (4/4)
gällande (6/6)
se (16/16)
noll (1/1)
relationsrådgivning (2/2)
km2 (5/5)
utsatt (23/23)
resekortet (2/2)
kostar (12/12)
ärekränkning (1/1)
handpenningen (1/1)
oavlönat (1/1)
skyldiga (4/4)
fackföreningsverksamhet (1/1)
skapar (1/1)
arbetskulturen (5/5)
rådgivningarna (2/2)
utlåtandet (3/3)
terminen (1/1)
uttrycka (2/2)
Nordea (1/1)
Kyrkbacken (1/1)
parktanterna (1/1)
preparaten (1/1)
banken (11/11)
diplomingenjörsexamen (1/1)
namn (21/21)
fritiden (1/1)
placera (2/2)
skadligt (1/1)
sök (1/1)
färdighetsnivå (2/2)
diskrimineras (6/6)
hjälpmedel (18/18)
punktlighet (3/3)
tidtabellerna (1/1)
konkurrenter (1/1)
ledd (5/5)
examina (8/8)
karriären (1/1)
skede (5/5)
konkurs (3/3)
räknare (1/1)
hemmaarbete (1/1)
skatterna (1/1)
ärende (3/3)
leta (7/7)
naturvetenskapliga (2/2)
varken (1/1)
boenderegistret (2/2)
övrigt (2/2)
stå (1/1)
utmätning (3/3)
undersida (1/1)
riksdagsval (2/2)
bostadsområde (4/4)
utvecklar (2/2)
individuella (1/1)
undervisnings- (1/1)
sända (1/1)
utländska (17/20) Utländska (3)
småbarnspedagogisk (1/1)
sådant (16/16)
lösa (2/2)
storleken (4/4)
arbetskontrakt (1/1)
hälsofrämjande (1/1)
API (1/1)
återvinning (6/6)
invandrararbetefinska (1/1)
CC (1/1)
problemen (1/1)
bekanta (6/6)
kollektivtrafikförbindelser (4/4)
historia (6/6)
grundundervisning (2/2)
yrkeshögskolor (9/12) Yrkeshögskolor (3)
Jourhjälpen (1/1)
Norden (1/1)
närmotion (1/1)
lokal (1/1)
betalar (71/71)
Luetaan (1/1)
jobbfinska (1/1)
istiden (1/1)
innehållet (4/7) Innehållet (3)
arbetat (10/10)
telefontjänst (11/11)
källskattekort (1/1)
ordna (23/23)
ungdomsarbetare (1/1)
gränsövergång (2/2)
stanna (10/10)
inlärnings- (1/1)
tider (10/10)
myndighetens (2/2)
surfplatta (1/1)
publiceras (1/1)
1500kt (1/1)
känna (6/6)
samlingar (3/3)
film (4/4)
Struves (1/1)
lokaltidningarna (1/1)
anhörig (9/9)
kyrkoherdeämbetet (1/1)
beteendefinska (3/3)
föräldraledighet (2/2)
ljusaste (1/1)
Furumo (3/3)
mångsidig (2/2)
upp (67/67)
organ (1/1)
fallen (1/1)
försäljningsmetoderna (1/1)
Nuorisoasuntoliitto (1/1)
änkling (2/2)
lähestymiskielto (1/1)
publicerades (1/1)
hautausavustus (1/1)
äktenskap (52/54) Äktenskap (2)
karriärmentorskap (1/1)
sexualitetfinska (1/1)
snöa (1/1)
instrument (2/2)
vapaaehtoisen (1/1)
vederbörligt (1/1)
bebott (3/3)
audiovisuella (1/1)
kilometer (2/2)
lönespecifikation (1/1)
jobbsajt (1/1)
inspiration (1/1)
ansiotulovähennys (1/1)
Europaskolan (1/1)
sjukdagpenning (11/11)
övernatta (5/5)
steg (5/5)
förmynderskap (2/2)
näringsbyråerfinska (1/1)
läskunnighet (1/1)
lösgjorde (1/1)
kommunens (18/18)
skeden (2/2)
yttre (1/1)
gränsöverskridande (1/1)
kompetensområden (1/1)
spis (1/1)
tidsfrist (2/2)
hitta (28/28)
hushållfinska (1/1)
socialmyndigheters (1/1)
kandidat (4/4)
Soite (5/5)
sexuell (5/5)
butiken (1/1)
packa (1/1)
vattenavgiften (3/3)
anslutningsblankett (1/1)
band (1/1)
Raumo (1/1)
gymnasieutbildning (6/6)
vita (4/4)
avkoppling (1/1)
förhindra (1/1)
hjälpsystem (1/1)
bankerna (1/1)
datoranvändningen (1/1)
lokala (8/8)
utvecklingsplan (2/2)
vinterlov (1/1)
enklast (1/1)
verk (1/1)
lekparkerna (1/1)
budskap (1/1)
koulukuraattori (1/1)
Facebook (1/1)
bor (84/84)
konkret (1/1)
sjukdomsfall (1/1)
samlar (1/1)
tidsbunden (2/2)
godkänd (3/3)
bioprogrammet (1/1)
hurudan (2/2)
Svartskär (1/1)
gränssnittet (1/1)
familjeärenden (2/2)
krig (4/4)
fasta (3/3)
avgörande (3/3)
upprättandet (3/3)
vänner (6/7) Vänner (1)
inleddes (2/2)
eftermiddagsverksamhet (3/3)
studielinjerna (1/1)
stödundervisning (3/3)
naturhuset (1/1)
ordningsnummer (1/1)
slidan (1/1)
konfidentiellt (3/3)
kuntoutustuki (1/1)
annons (1/1)
sorgfinska (1/1)
röst (3/3)
grundlagen (2/2)
samhället (14/14)
valkretsen (1/1)
gifte (1/1)
dagvårdfinska (3/3)
sämre (3/3)
bankkonto (14/14)
käsiraha (1/1)
webbplatserna (1/1)
volontärarbetefinska (1/1)
åldrarna (2/2)
pedagoger (2/2)
komihåglista (2/4) Komihåglista (2)
företagsrådgivningscentra (1/1)
huvudhälsostationen (1/1)
bedömningsgrunder (1/1)
linor (1/1)
inget (21/21)
upptäckande (1/1)
palveluohjaaja (1/1)
parterapi (1/1)
vad (22/24) Vad (2)
långvarig (3/3)
markägarna (1/1)
heltid (8/8)
motionsspår (1/1)
svagheterna (1/1)
Firmaxifinska (1/1)
försörjningen (4/4)
skattebyråns (1/1)
kartläggs (1/1)
stadsdelfinska (3/3)
näringsbyrån (40/40)
korkein (1/1)
Bredvikens (1/1)
Sporttikortti (1/1)
väsentlig (3/3)
fortlöpande (2/2)
goda (10/10)
Verla (1/1)
siktar (1/1)
mödrahem (2/2)
utsökningfinska (1/1)
besegrat (1/1)
köpte (1/1)
ändrade (1/1)
tvåspråkigt (2/2)
presidentvalfinska (1/1)
kansainvälinen (1/1)
beror (42/42)
folk (2/2)
bedömning (6/6)
Nödcentralsverkets (1/1)
fisk (1/1)
länderfinska (1/1)
andelslagets (3/3)
biojäte (1/1)
handikapp (18/18)
upprätta (6/6)
lägga (5/5)
hyresvärder (1/1)
europeiska (11/18) Europeiska (7)
relationer (1/1)
tekniska (1/1)
religionssamfund (4/4)
lekpark (2/2)
onsdag (1/1)
väcker (3/3)
kortet (8/8)
högskolexamenfinska (1/1)
befriats (2/2)
vägguttaget (1/1)
erkännande (12/14) Erkännande (2)
föra (12/12)
järnvägsstationer (1/1)
jobbförmedlingssidor (2/2)
detaljerna (1/1)
ingriper (1/1)
reglerade (4/4)
arbetarskyddsmyndigheternafinska (1/1)
amatörteatrar (2/2)
Halloween (1/1)
dans (6/6)
bostäder (38/38)
työttömyysturvan (1/1)
anställd (15/15)
innehavarkort (1/1)
motionstjänsternafinska (1/1)
erkänns (1/1)
alltför (3/3)
post (32/32)
reseförsäkring (1/1)
anpassa (1/1)
Tysklands (1/1)
gåvor (1/1)
skatteräknare (1/1)
päivystys (3/3)
existerande (1/1)
elarbeten (1/1)
gravområde (2/2)
redaktioner (1/1)
kris (2/2)
sukupuolitauti (1/1)
min (5/7) Min (2)
Tullens (1/2) tullens (1)
visumcentralen (1/1)
sortering (1/1)
ifrån (5/5)
alls (1/1)
sällskapar (1/1)
rådgivningen (23/23)
tillväxten (1/1)
församlingar (10/10)
moderna (1/1)
friska (1/1)
initiala (2/2)
brotten (1/1)
producera (3/3)
rådgivningsbyråernas (2/2)
hyresbostaden (2/2)
80:e (1/1)
mental- (2/2)
uteblir (1/1)
Hagalunds (1/1)
måsta (1/1)
vuxenläroanstalter (2/2)
rösträtt (13/13)
Pyhäjoki (1/1)
uppgifter (37/39) Uppgifter (2)
familjepensionen (1/1)
räddningsverk (1/1)
turistbyrå (1/1)
hyresgästerna (1/1)
avgår (2/2)
egenskaper (1/1)
parkeringsbiljetten (1/1)
majoriteten (1/1)
polikliniken (8/8)
hörselskadade (5/5)
naken (1/1)
pensionerad (1/1)
Nelonen (1/1)
hälsopunkterfinska (1/1)
hoppas (1/1)
minuter (1/1)
privatvårdsstödet (1/1)
rakt (3/3)
läs (2/2)
svår (5/5)
kran (1/1)
Nationalgalleriet (1/1)
boende (44/48) Boende (4)
färger (1/1)
dispens (2/2)
kuljetuspalvelu (1/1)
medborgarskapsansökan (2/2)
utbildnings (1/1)
studieförmåga (1/1)
befolkningen (3/3)
sortera (1/1)
ägaren (1/1)
minipiller (1/1)
Monikas (1/1)
söderifrån (1/1)
förlossningsavdelning (1/1)
arbetslöshetspenning (1/1)
karta (1/1)
koulu- (1/1)
lokaler (7/7)
servicecentret (1/1)
erkänts (3/3)
liv (15/15)
registrerad (3/3)
Mannerheims (2/2)
öppna (55/55)
orsakar (4/4)
landskapsbibliotek (3/3)
terveysministeriö (2/2)
alkohol (6/6)
inkluderar (1/1)
vägar (1/1)
tillverkas (2/2)
bistår (2/2)
vuxenutbildningen (1/1)
kulturkontor (1/1)
bussar (4/4)
vaccinationsprogrammet (1/1)
arbetslöshetskassafinska (1/1)
lämpar (2/2)
elevens (8/8)
smärtor (3/3)
hembygdsmuseerna (1/1)
samt (81/81)
undervisas (3/3)
specialgymnasier (1/1)
höjs (1/1)
arbetslöshetsförsäkringen (2/2)
idrottsplatser (5/5)
duar (3/3)
planen (1/1)
ansvarig (4/4)
utvisas (2/2)
tagit (2/2)
företagarhandböcker (1/1)
övertygelse (5/5)
handlingar (11/11)
Registreringsanmälan (1/2) registreringsanmälan (1)
EES (35/35)
bosättningsbaserade (1/1)
tullanmäla (1/1)
kontonummerfinska (1/1)
ägare (6/6)
England (1/1)
garanterar (1/1)
hyresgästenfinska (1/1)
nummer (6/6)
läkarens (2/2)
tutkiminen (2/2)
resmål (1/1)
slutligen (1/1)
kyrkanfinska (1/1)
beskickningar (10/10)
lagenliga (1/1)
åtta (3/3)
stugan (1/1)
pensionsanstalt (3/3)
myndigheter (35/35)
ungdomars (1/1)
trafiken (2/3) Trafiken (1)
speciellt (9/9)
bestämd (4/4)
riskerna (1/1)
nödvändiga (5/5)
utvecklas (2/2)
tjänstemännen (2/2)
repetera (1/1)
Närpes (1/1)
temadagar (1/1)
preventivrådgivning (1/1)
turist (2/2)
lånas (1/1)
hobbyutbud (1/1)
förskolebarn (2/2)
bilhandlare (1/1)
skrivna (1/1)
vattenkonsumtionen (1/1)
framstegsvänligt (1/1)
som (1265/1266) Som (1)
returnera (1/1)
anges (11/11)
högtid (1/1)
kapitalinkomst (1/1)
mångfald (2/2)
medan (5/5)
återhämta (2/2)
hyresvärdens (2/2)
godkänts (3/3)
växelvis (1/1)
samiska (8/8)
fackliga (1/1)
instruktioner (1/1)
terveysasema (13/13)
startandet (1/1)
grundar (6/6)
stödengelska (1/1)
arbetsintervju (1/1)
byrå (17/17)
vistas (35/35)
ombord (1/1)
perustuslaki (1/1)
bilskola (1/1)
folkhögskolafinska (1/1)
konserter (1/1)
licensen (2/2)
socialstationen (1/1)
arvolautakunta (1/1)
fyllas (1/1)
garantipensionen (2/2)
allmänheten (2/2)
sådan (9/9)
alternativen (1/1)
knöt (1/1)
tungt (1/1)
dyra (6/6)
anslagstavlor (1/1)
autonoma (1/1)
eventuell (2/2)
övrig (2/2)
fallet (2/2)
religion (31/31)
kulturcenter (1/1)
överföras (1/1)
anhörigafinska (1/1)
anställa (3/3)
arbetsplats (27/27)
nationer (1/1)
företaget (18/18)
städernas (1/1)
pensionärerfinska (1/1)
-årigt (1/1)
rådgivningstjänst (5/5)
skedet (1/1)
musicera (1/1)
sagts (1/1)
kundtjänstfinska (1/1)
prioriteras (2/2)
stödet (12/12)
bör (18/18)
tomt (1/1)
väg (2/2)
tvingade (1/1)
kemikaler (1/1)
borgare (1/1)
yrkesbevis (1/1)
utlandsprefix (1/1)
bakgrundsmusik (2/2)
gymnasieskolorna (2/2)
klarspråk (1/1)
skuldfria (1/1)
hemfrid (1/1)
arbetssökanden (1/1)
sägas (2/2)
ras (2/2)
bibehålls (1/1)
Marthaförbundetfinska (1/1)
arbetsavtal (8/8)
arbetspensionsutdragen (1/1)
välfärds- (1/1)
Arctica (3/3)
busstation (1/1)
asumisoikeussopimus (1/1)
rusmedelsberoende (1/1)
teoretiska (1/1)
dagpenning (13/13)
ålderspensionsålder (1/1)
gånger (13/13)
vädra (1/1)
kostnadsfria (11/11)
träffa (8/8)
mor (11/11)
köpet (4/4)
flyktingfinska (1/1)
specialdiet (1/1)
joustava (1/1)
pensionsanstalten (1/1)
Menyn (1/2) menyn (1)
kontakt (51/51)
nämnda (3/3)
gruppmöten (1/1)
konsumtionsskatt (1/1)
förtroendeman (4/4)
uppvisa (1/1)
harmoniska (1/1)
drivs (5/5)
familjeåterförening (6/6)
hittat (3/3)
överklaga (7/7)
rehabiliteringsstöd (1/1)
flygplatsen (1/1)
rekisteröintitodistus (2/2)
flyttningen (3/3)
nätetfinska (1/1)
fuktproblem (1/1)
övriga (28/28)
språketfinska (6/6)
-svenska (1/1)
råkat (4/4)
missbruks- (1/1)
leker (1/1)
sjukhusavgifter (1/1)
textfält (1/1)
egenvårdsläkemedel (1/1)
information (337/342) Information (5)
magisterexamen (3/3)
domstol (2/2)
sådana (14/14)
tillsvidare (6/6)
vuxenutbildning (8/8)
slutfört (1/1)
tolka (1/1)
rekommendabelt (1/1)
varannan (1/1)
meddelande (4/4)
asuntosäätiö (2/2)
gottgörelse (1/1)
underteckna (4/4)
hälstocentralen (1/1)
fler (10/10)
grädde (1/1)
legitimerad (1/1)
stavelsen (1/1)
invandrafamiljer (1/1)
sökmotor (6/6)
dagen (15/15)
läroboken (1/1)
omgivningen (1/1)
småbarnspedagogiken (12/12)
strykjärnet (1/1)
socken (1/1)
anordnar (1/1)
Kuluttajansuojalaki (1/1)
identiska (3/3)
dagvårdsplatserfinska (1/1)
HSL (2/2)
bensinstationer (2/2)
kostnaderna (15/15)
återhämtar (3/3)
bostadsförsäljningsannonser (2/2)
beslutsmakt (1/1)
begränsat (1/1)
beräknas (10/10)
borta (1/1)
filmarkiv (1/1)
ansökningarna (2/2)
västländerna (1/1)
sökande (6/6)
sorggrupper (1/1)
Mielenterveys (1/1)
punktligt (1/1)
hammashoito (1/1)
nödläge (1/1)
finansierat (1/1)
progressiv (4/4)
trots (6/6)
krigen (2/2)
hemkommun (104/114) Hemkommun (10)
läkemedelfinska (1/1)
stambyte (1/1)
övningar (1/1)
arbetsmarknaden (1/1)
hit (1/1)
magistratet (1/1)
kieli (1/1)
grundlag (2/2)
valkrets (1/1)
identiteten (2/2)
konst (11/12) Konst (1)
läroverket (1/1)
beaktande (2/2)
statliga (9/9)
storlekar (1/1)
köpt (3/3)
minderårigt (4/4)
femte (2/2)
hälsovårdenfinska (1/1)
förälderns (3/3)
landsomfattande (1/1)
thai (10/10)
ägs (9/9)
kommunikationsfärdigheter (1/1)
neutral (1/1)
semester (4/4)
specialvårdspenning (1/1)
betalningsanmärkningar (2/2)
viseringsfria (1/1)
födelsedatum (3/3)
hälsovårdscentraler (1/1)
platsansökan (1/1)
kulturarvet (1/1)
vårdnaden (8/8)
rösten (1/1)
intyg (26/26)
inleds (8/8)
fönstren (2/2)
fiske (3/3)
personbolag (1/1)
3D (1/1)
makars (1/1)
arbetarskyddfinska (2/2)
Trafi (1/1)
Sparbanken (1/1)
grunda (31/31)
tidsbegränsade (1/1)
oppisopimustoimisto (1/1)
längd (3/3)
säkert (3/3)
minnesbilderna (1/1)
helhet (3/3)
regelbundet (5/5)
gift (12/12)
folkhögskolan (3/3)
förlossning (8/8)
webbtjänst (9/9)
tuberkulosfinska (2/2)
möter (1/1)
teoretiskt (1/1)
uppfylla (3/3)
huvudansvaret (1/1)
behåller (2/2)
oman (1/1)
gårdsbyggnader (1/1)
heller (14/14)
riksomfattande (4/4)
utvecklingsstörd (3/3)
registreringen (6/6)
ländernafinska (1/1)
kommunalval (9/9)
interna (1/1)
fråga (68/68)
webbundervisning (1/1)
ökat (3/3)
militärunderstöd (1/1)
överklagar (1/1)
utfärdades (1/1)
olycksfallsförsäkring (3/3)
dagvårdens (2/2)
satt (2/2)
påminnelse- (1/1)
inverka (1/1)
ungdomscentralen (1/1)
utnyttjande (1/1)
underlivet (1/1)
idka (4/4)
posten (2/2)
marker (1/1)
delvis (10/10)
kb (4/5) kB (1)
Global (7/7)
år (260/260)
diabetesfinska (1/1)
upphovsrätts- (1/1)
brister (3/3)
VR:s (2/2)
arbetstider (5/5)
vårdåtgärder (1/1)
barnuppfostran (1/1)
inloggning (1/1)
exempelvis (15/15)
ålderspensionen (3/3)
äldrefinska (1/1)
intyga (1/1)
vitsorden (1/1)
svar (1/1)
politik (1/1)
tillåtet (6/6)
senaste (9/9)
träffar (1/1)
rädd (3/3)
publicus (2/2)
företagsformen (3/3)
grund (122/122)
påtryckningar (1/1)
motionsevenemang (1/1)
primärhälsovård (2/2)
informationsförmedlare (1/1)
tidsbegränsat (2/2)
studieområden (4/4)
krävande (5/5)
tolkcentraler (2/2)
betalt (2/2)
tjänstestyrningen (1/1)
varmare (1/1)
magisterstudierna (1/1)
startpenningen (1/1)
näringsministeriet (8/8)
husbolagets (2/2)
Företagsrådgivning (2/4) företagsrådgivning (2)
producerar (1/1)
arbetstagarnas (5/5)
högskolorna (7/7)
polikliniker (2/2)
språkcaféer (2/2)
ekonominfinska (1/1)
nödvändigt (4/4)
socialverk (2/2)
orsaka (5/5)
sina (57/57)
förbjudet (2/2)
rättshjälpen (1/1)
pojkar (4/4)
Institutet (2/3) institutet (1)
urspråken (1/1)
speciella (1/1)
folkhögskolorfinska (1/1)
småstad (1/1)
idrottsmöjligheter (2/2)
arbetslandet (1/1)
erövrades (1/1)
sjuk- (1/1)
namnen (3/3)
bank (4/5) Bank (1)
Helsingforstilläggetfinska (1/1)
suomi.fi (2/3) Suomi.fi (1)
panelen (2/2)
utvecklingsidéer (1/1)
gatan (1/1)
dagvårdsproducenten (1/1)
föräldrarnafinska (1/1)
symtom (1/1)
arbetslös (34/34)
skyddshem (15/18) Skyddshem (3)
kostnad (1/1)
webben (2/2)
fortbildar (1/1)
vattendrag (3/3)
sökmotorer (1/1)
snabba (1/1)
servicevägledning (1/1)
doula (1/1)
studieplaner (1/1)
legaliserat (2/2)
räkning (3/3)
bankgiroblankett (1/1)
Clinic (7/7)
granne (6/6)
heder (1/1)
slutsyn (1/1)
preparat (1/1)
restaurangbranschen (1/1)
driver (3/3)
näringar (1/1)
familjeförhållande (1/1)
vårdens (1/1)
livsåskådningskunskap (2/2)
biblioteks (1/1)
möjligheterna (3/3)
finns (411/411)
understiger (1/1)
medborgarna (2/2)
ombes (1/1)
ammattiliitto (1/1)
bibliotekskunderna (1/1)
annanstans (10/10)
webbläsarinställningar (1/1)
besöken (1/1)
läkarstationfinska (1/1)
idrottshobbyer (1/1)
utrikesflygen (1/1)
tandvårdsjouren (1/1)
religioner (3/4) Religioner (1)
handikapptjänster (2/2)
anställningstiden (1/1)
fall (62/62)
grammatikfinska (1/1)
baserar (1/1)
bolsjevikregeringen (1/1)
kunnat (2/2)
Rysslands (2/2)
lönebesked (1/1)
arbetet (49/49)
orsak (7/7)
inkludera (1/1)
studentexpeditionen (1/1)
effektiva (1/1)
lagstadgad (2/2)
kiinteistövero (1/1)
yrkesutbildningenfinska (1/1)
tågen (1/1)
opintotuki (2/2)
nyttar (1/1)
arbetsvillkoret (2/2)
kontanter (5/5)
programmeringsgränssnitt (1/1)
universitetets (2/2)
teatrar (4/4)
hög (7/7)
distansstudier (1/1)
osittainen (1/1)
kurdiska (24/24)
socialt (1/1)
yrkeskvalifikationer (1/1)
promenader (1/1)
C2 (1/1)
församlingarna (4/4)
förlossningsdatum (1/1)
landsbygden (3/3)
semesterersättning (2/2)
blev (17/17)
Nivavaara (1/1)
funktionshinder (1/1)
underhållsskyldiga (1/1)
tänkande (1/1)
viseringspliktigt (1/1)
förvalta (2/2)
barntillsynsmannen (1/1)
hitar (2/2)
gångtrafiken (1/1)
resenärerfinska (1/1)
avtog (1/1)
hoitotakuu (1/1)
våningen (4/4)
finansieringsalternativ (3/3)
bassjälvrisk (1/1)
underskrifterna (1/1)
männen (1/1)
snabb (1/1)
moderskaps- (1/1)
Työväen (2/2)
motionärer (1/1)
lätt (5/5)
barnrådgivningen (8/8)
originalspråk (1/1)
köparens (1/1)
stegen (1/1)
nätverka (1/1)
kontrollera (19/19)
avlidnes (2/2)
stöd (81/92) Stöd (11)
väster (2/2)
lägsta (1/1)
rättsväsendet (1/1)
sjukfall (3/3)
hälsomotionskalendern (1/1)
bytet (1/1)
Kärlek (1/1)
företagsformer (2/3) Företagsformer (1)
burmesiska (1/1)
Mejlansvägen (1/1)
biljettkontoren (1/1)
spisen (4/4)
gardinerna (1/1)
delges (1/1)
fortbildningfinska (1/1)
inkvartering (2/2)
vähennykset (1/1)
produktionen (1/1)
närvarande (3/3)
kommunicerar (1/1)
polisanmäla (1/1)
telefonjouren (1/1)
varmaste (1/1)
akuta (5/5)
jobbsajter (2/2)
skuldrådgivning (3/3)
julgran (1/1)
förvärvsinkomstavdrag (1/1)
insjöarna (1/1)
sälj (1/1)
trafikverkets (1/1)
semesterresor (1/1)
torra (2/2)
universitetssjukhus (2/2)
servicecenter (1/1)
översättningarna (1/1)
uttryckligen (1/1)
kundens (2/2)
återkallande (1/1)
stunder (1/1)
handledd (2/2)
originalspråket (1/1)
lagen (26/26)
europeiskt (2/2)
verket (9/9)
somliga (1/1)
träning (1/1)
vårdas (8/8)
påverkan (5/5)
romanifinska (1/1)
sjukvårdfinska (1/1)
religionen (2/2)
hurdan (2/2)
anstalt (2/2)
samhällsvetenskaper (2/2)
praktik (4/4)
beslut (47/47)
statsstöd (1/1)
samtycke (4/4)
nätter (1/1)
helger (6/6)
rådfråga (2/2)
nia (2/2)
föräldraledigheten (7/7)
äktenskapsintyg (4/4)
ändringar (6/6)
cykling (4/4)
simpass (1/1)
företagshälsovårdens (1/1)
ämnet (6/6)
bygga (6/6)
miljöministeriet (1/1)
registerstyrelsens (1/1)
kandidater (1/1)
avliden (1/1)
statsministern (2/2)
distansgymnasiet (1/1)
insulin (1/1)
anarki (2/2)
tre (83/83)
sakkunskap (1/1)
arbetslöshetsersättning (10/10)
studielinjer (1/1)
vuxengymnasiums (1/1)
grundläggande (43/45) Grundläggande (2)
hobbyredskap (1/1)
specialboende (1/1)
rosoll (1/1)
ungdom (1/1)
tilläggsutbildning (3/3)
kunnanvaltuusto (1/1)
små (15/15)
inför (11/11)
finlandssvenskarna (1/1)
ihop (1/1)
byggdes (1/1)
månaden (6/6)
inskärper (1/1)
tillståndsansökan (4/4)
danskonst (1/1)
angelägenheter (5/5)
snabbt (11/11)
namnet (2/2)
varhaiskasvatushakemus (1/1)
kommunfullmäktige (5/5)
beskickningen (14/14)
byar (1/1)
anstaltsvårdenfinska (1/1)
anonymt (2/2)
viktig (15/15)
apotekets (3/3)
B (7/7)
studerandena (1/1)
följas (1/1)
oktober (2/2)
löpt (2/2)
bosatt (19/19)
hänvisa (1/1)
Ristin (2/2)
presenter (2/2)
köptjänst (1/1)
terminsavgifter (1/1)
delarna (2/2)
jämlikt (4/4)
plågor (1/1)
byråerna (1/1)
lyfta (3/3)
språk- (3/3)
makthavaren (1/1)
barnskyddet (4/4)
hjälpbehovet (2/2)
föregår (1/1)
Tammerforsregionen (1/1)
hälsoproblem (1/1)
lagakraftvunnet (1/1)
hemhjälp (1/1)
idrottssällskap (2/2)
utevistelser (2/2)
skattedeklaration (1/1)
utbetalad (2/2)
upphovsrättsliga (1/1)
föreslår (3/3)
kunna (38/38)
asylprocessen (1/1)
grannmedling (1/1)
ses (1/1)
omhändertas (1/1)
järnvägsstationerna (1/1)
gruppera (1/1)
lastensairaala (1/1)
språkanvändares (2/2)
viseringsskyldiga (1/1)
vilkas (1/1)
utflykter (6/6)
grunder (9/9)
yrkesbeteckning (1/1)
ställs (5/5)
konstindustri (2/2)
tatarer (1/1)
säker (5/5)
medeltida (1/1)
helgons (3/3)
työ- (3/4) Työ- (1)
sig (184/184)
kort (21/22) Kort (1)
betala (88/88)
enskilda (6/6)
fisket (1/1)
bostadfinska (3/3)
semesterdagar (1/1)
tack (4/4)
stannar (5/5)
användningen (6/6)
Barnsjukhuset (2/3) barnsjukhuset (1)
pensionssystem (1/1)
A1.1 (1/1)
beslutat (2/2)
ingendera (1/1)
kollektivavtalen (3/3)
enlighet (7/7)
parförhållandet (14/14)
konstskola (1/1)
julstjärnor (1/1)
krisen (1/1)
kunskap (2/2)
Nyland (8/8)
beslutas (5/5)
bekänna (1/1)
asylansökan (15/15)
arbetsoförmögenhet (2/2)
läkemedlet (3/3)
440kt (1/1)
at (3/3)
Apostille (1/1)
anspråkslös (1/1)
hemförsäkringen (4/4)
perioder (5/5)
barnskyddsmyndigheten (2/2)
högklassig (1/1)
församlingssammansutning (1/1)
Europa (3/3)
fostras (2/2)
skuldrådgivningen (1/1)
växlande (1/1)
VAV (2/2)
avträdelseanmälan (1/1)
osakliga (1/1)
bäst (9/9)
grundexamen (7/7)
typ (4/4)
veronumero (2/2)
punkt (1/1)
röra (20/20)
emot (13/13)
trakasserar (1/1)
gymnasieskolans (1/1)
Tyttöjen (1/1)
åtföljs (2/2)
vigselförrättningen (1/1)
papperslösa (6/6)
stadssund (1/1)
rädsla (1/1)
mammor (1/1)
juridik (2/2)
identifierats (1/1)
centraliserade (3/3)
tillväxt (4/4)
toimintakeskus (1/1)
handikappade (35/36) Handikappade (1)
Koivuhaan (1/1)
arbetsmarknadsstödets (1/1)
vägande (5/5)
elva (3/3)
skyddsbehov (1/1)
hoitoraha (2/2)
överklagan (1/1)
tills (16/16)
kranen (1/1)
begravningen (3/3)
möjligtvis (1/1)
utländskt (2/2)
Vinge (2/2)
ventilationssystem (1/1)
skapade (1/1)
jaga (1/1)
plan (1/1)
flytten (7/7)
studentkår (1/1)
grundskolor (4/4)
familjehus (1/1)
arvingarna (1/1)
arbetstagarens (5/5)
kulturen (10/10)
sysselsättning (5/5)
orsaker (8/8)
evangelisk (17/17)
hemvist (2/2)
funktionellt (1/1)
flyktinghjälp (3/3)
nedsättande (2/2)
gruppfamiljedagvården (1/1)
fett (1/1)
asumisoikeusmaksu (1/1)
Karlebynejden (1/1)
Myyringin (1/1)
respons (6/6)
fakturera (2/2)
firas (11/11)
organisera (1/1)
församlingen (1/1)
avsätta (1/1)
köa (1/1)
kriget (4/4)
anor (1/1)
arbetsmarknadsstödet (1/1)
socialservicecenter (1/1)
föreskriver (1/1)
förtroende (1/1)
modersmålet (6/6)
besvara (1/1)
lugga (1/1)
tvungen (8/8)
förknippas (1/1)
Uudenmaan (1/1)
hel (1/1)
åka (5/5)
kulturstad (1/1)
ansökningstiderna (2/2)
ort (5/5)
Renlund (1/1)
boka (57/57)
bådas (2/2)
övernattar (1/1)
familjeplaneringfinska (2/2)
ingår (23/23)
spänning (2/2)
A1 (5/5)
opetus (2/2)
teaterfinska (1/1)
synskadades (1/1)
västeuropéer (1/1)
förarutbildning (1/1)
grannar (1/1)
skadad (1/1)
fostret (1/1)
förvänta (1/1)
nödsituationer (8/8)
picknick (1/1)
stödundervisningen (1/1)
lönerna (3/3)
asiointi (1/1)
fisketillstånd (3/3)
herpes (1/1)
avses (16/16)
privatpersoner (8/8)
uppehållstillståndfinska (6/6)
utbildningskoncern (1/1)
verksamhetssätt (1/1)
haltijakohtainen (1/1)
kämpade (1/1)
maahanmuuttajapalvelut (1/1)
rådgivningstjänster (4/4)
grundskola (1/1)
centraliserat (1/1)
oleskeluoikeuden (1/1)
praktikant (1/1)
närheten (4/4)
gravkontor (1/1)
böter (4/4)
elektroniska (5/5)
motiverat (1/1)
rättshjälp (5/5)
översättningen (4/4)
största (16/16)
miljöcentralerna (1/1)
egnahemshus (5/5)
missbrukat (1/1)
ledigheten (1/1)
skild (1/1)
Informationscentralen (2/2)
brottsoffret (1/1)
fram (13/13)
frukta (1/1)
utsänd (1/1)
haft (7/7)
övervåningen (1/1)
unionenfinska (1/1)
löntagar- (1/1)
nattcaféet (1/1)
telefon (38/38)
bekostat (1/1)
tandhälsovårdenfinska (1/1)
rådgivningsbyråns (1/1)
öppettider (8/8)
arbetsinkomster (2/2)
tillgång (5/5)
vårdartiklar (1/1)
kring (9/9)
Sandudd (1/1)
bekostas (1/1)
helgerna (2/2)
förbjuder (5/5)
flyttningsdagen (1/1)
nätterna (3/3)
elapparat (2/2)
landskommunen (1/1)
hoitoapupalvelu (1/1)
elden (1/1)
umgängesrättfinska (2/2)
inrättas (1/1)
äkta (1/2) Äkta (1)
transport (1/1)
volym (1/1)
fyrverkerier (1/1)
fastställas (3/3)
daghemfinska (1/1)
makans (1/1)
förfaller (2/2)
valmistava (1/1)
Eira (1/1)
oktoberrevolutionen (1/1)
företagets (8/8)
kl. (1/1)
bostadslånet (3/3)
kielenkäyttäjän (2/2)
kuntoutuspsykoterapia (1/1)
vin (1/1)
ändra (6/6)
räntan (2/3) Räntan (1)
vart (10/10)
flyttades (2/2)
valtion (1/1)
Bio (1/1)
vaginalt (2/2)
förteckning (5/5)
arbetspensionsutdraget (1/1)
överklagas (1/1)
insinööri (1/1)
frivilligarbeta (1/1)
styrkor (1/1)
inkomstgränsen (1/1)
ruokakunta (1/1)
Asokoditfinska (2/2)
prövningfinska (2/2)
virkatodistus (1/1)
betraktar (1/1)
Kylämaja (1/1)
Helsingforsregionens (10/10)
siviilisäätytodistus (1/1)
fel (12/12)
stöds (1/1)
ränta (1/1)
fick (12/12)
arbetafinska (2/2)
specialkompetens (1/1)
ArPL (1/1)
möten (6/6)
höst (1/1)
FPA.I (1/1)
skilda (1/1)
fastighet (4/4)
noggrant (2/2)
tecknat (1/1)
tillrådligt (1/1)
byråer (3/3)
skolkuratorerna (2/2)
pysyvä (1/1)
bostadsansökan (3/3)
invandrarbakgrund (5/5)
social- (26/26)
giltighetstid (1/1)
hemort (17/17)
underhållsförmåga (2/2)
situation (31/31)
läget (1/1)
värnpliktiga (1/1)
stipendiesystem (2/2)
erbjuda (3/3)
omskärelse (6/6)
rektorn (1/1)
skolgång (4/4)
tvingats (1/1)
följebrev (1/1)
barnbidrag (8/9) Barnbidrag (1)
gång (14/14)
konstmuseum (2/2)
webbplatsens (1/1)
språkkunniga (1/1)
prov (6/6)
drar (1/1)
körkort (11/11)
normalt (4/4)
mångkulturellt (2/2)
magistratens (7/7)
Clubs (1/1)
grunddagpenning (8/8)
nyttigt (2/2)
försörjning (12/12)
sektorn (10/10)
smal (1/1)
tillståndskort (1/1)
Rovaniemifinska (2/2)
Island (7/7)
Soldatskär (1/1)
måltid (2/2)
International (2/2)
turvapaikkapuhuttelu (1/1)
säkring (1/1)
evenemangskalendrarna (3/3)
ägarbostäder (1/1)
funktionsförmåga (1/1)
sosiaalitoimisto (3/3)
Project (1/1)
ungdomsledarna (1/1)
tolv (6/6)
representerade (4/4)
läkarpriserfinska (1/1)
framskrider (3/3)
kännedom (1/1)
affärsverksamheten (2/2)
flyttas (1/1)
midnattssolens (1/1)
etniska (3/3)
hyresgäster (3/3)
förändrades (1/1)
syskonrabatt (1/1)
tillräcklig (10/10)
Hakunilan (1/1)
halvsyskon (1/1)
privatvårdsstöd (2/2)
uppståndelse (1/1)
status (1/1)
grundande (3/3)
måndag (9/9)
begränsar (2/2)
utredningar (5/5)
familjeplaneringsrådgivningarna (1/1)
påtryckning (1/1)
gott (7/7)
sysselsättningstjänster (1/1)
Oikarainen (1/1)
skorna (1/1)
www.teosto.fi (1/1)
söks (4/4)
lågstadiets (1/1)
sluttexterna (1/1)
avtalet (21/21)
jämställdhetsombudsmannen (3/3)
Centralorganisation (1/1)
sigfinska (1/1)
registerstyrelsen (5/5)
disponent (2/2)
uppförande (1/1)
makarna (18/18)
giltigt (12/12)
stängda (2/2)
klockan (10/10)
vägg (1/1)
betalningsstörningfinska (1/1)
prat (2/2)
experter (3/3)
bakgrund (5/5)
kejsarsnitt (3/3)
pass (23/23)
yrkessjukdom (1/1)
egen (83/83)
beakta (7/7)
tandvårdsjourenfinska (1/1)
kommunal (6/6)
prövotiden (2/2)
korttidsvård (1/1)
psykiatriskötare (1/1)
uppförs (1/1)
avboka (2/2)
anskaffningspris (1/1)
mentalvårdstjänsterna (1/1)
tulosyksikkö (1/1)
koulukuraattorit (1/1)
tandläkarkontroller (1/1)
meriterna (1/1)
förening (9/9)
föräldrapenning (3/3)
hälsoåvård (1/1)
inkomstbeskattningfinska (1/1)
skattepengarna (1/1)
utlänningar (19/19)
ner (4/4)
säsongsarbetsvisum (1/1)
skiftarbetstillägg (1/1)
ordnade (1/1)
broschyren (1/1)
studiepenning (2/2)
tigga (1/1)
lönekvittona (1/1)
badar (4/4)
MERCURIA (1/1)
dragits (1/1)
partner (12/12)
förmedlar (2/2)
Förbundfinska (1/1)
svars (1/1)
parförhållandets (1/1)
yhdenvertaisuuslaki (1/2) Yhdenvertaisuuslaki (1)
reda (22/22)
flaskor (1/1)
tyger (1/1)
grunddagpenningen (1/1)
delat (1/1)
familjedagvård (2/2)
tillverka (1/1)
närskola (3/3)
klinikkaan (1/1)
avtalas (1/1)
stadigt (1/1)
överförda (1/1)
gränser (2/2)
receptbelagda (1/1)
existerar (3/3)
kamratstöd (2/2)
Skatteförvaltningens (9/12) skatteförvaltningens (3)
webbtjänsten (7/7)
egenföretagare (1/1)
kriser (1/1)
godkänner (4/4)
beskrivningar (1/1)
äidinkielen (1/1)
Konsumentförbund (1/1)
psykologi (1/1)
Trapesa (2/2)
idkas (2/2)
kartlägga (2/2)
inhyste (1/1)
sakkunnig (2/2)
författningar (1/1)
förverkligandet (1/1)
nycklarna (1/1)
tandvårdstjänsterna (1/1)
tävlingsdeltagaren (1/1)
ökade (1/1)
Kuntien (1/1)
tvunget (1/1)
pensionskassor (2/2)
myndigheterna (16/16)
pappfabrik (1/1)
vuxensocialarbetet (1/1)
Rinteenkulmafinska (1/1)
tredje (6/6)
gardena (1/1)
gårdar (1/1)
gymnasiernas (1/1)
förekomma (2/2)
åstadkomma (1/1)
klädskåp (1/1)
olägenhet (1/1)
anställningsvillkor (1/1)
hända (2/2)
kaupunki (1/1)
ordföranden (3/3)
Rovala (2/2)
kalendern (1/1)
narkos (1/1)
politisk (2/2)
hyresstöd (2/2)
till (1547/1553) Till (6)
frivilligt (8/8)
efter (88/88)
samerna (1/1)
gymnasium (13/14) Gymnasium (1)
upplevt (1/1)
varderas (1/1)
satsat (1/1)
meddelandekortet (1/1)
sjukdom (20/20)
informationen (6/6)
kamratförening (1/1)
ortodoksinen (1/1)
skattenummer (5/5)
studier (80/81) Studier (1)
servicesställen (1/1)
yrkeshögskolorfinska (4/4)
verksamhetsställe (6/6)
larmar (1/1)
världskriget (2/2)
dagvårdsenhet (1/1)
College (1/1)
glömde (1/1)
betraktas (5/5)
ljus (2/2)
ändå (25/25)
samjouren (1/1)
företagare (51/54) Företagare (3)
tillhandahållas (1/1)
sträckte (1/1)
digital (1/1)
nätet (13/13)
användning (2/2)
bildas (4/4)
lånegaranti (1/1)
få (338/338)
långfredagen (1/1)
Kokkola (2/2)
också (308/308)
äventyras (1/1)
avoin (7/7)
läs- (1/1)
myndighetshandlingen (1/1)
broschyrer (2/2)
svenskspråkigt (4/4)
arbetssökandefinska (2/2)
lager (1/1)
fullmäktiges (2/2)
marken (1/1)
belägen (1/1)
tillfällig (9/9)
familjerfinska (3/3)
åtalsprövning (1/1)
ekonomi (4/4)
kondition (1/1)
finansierar (1/1)
Akademi (1/1)
disponibla (3/3)
A1.2 (1/1)
Pro (3/3)
teaterfestivaler (1/1)
Europaparlamentet (4/4)
föreningsmötet (1/1)
andra (185/185)
ordningen (1/1)
verohallinto (1/1)
tis (2/2)
oppisopimuskoulutus (1/1)
webbplatser (13/13)
erhöll (1/1)
bulgariska (6/6)
ställning (9/9)
desto (1/1)
Konttisen (1/1)
arbetsplatserna (7/7)
salar (1/1)
juridisk (7/7)
Anon (1/1)
rekryteringsevenemang (1/1)
viga (1/1)
avoimet (2/2)
affärsverksamhetsplan (9/9)
religiöst (9/9)
medgivande (3/3)
mopedkort (1/1)
r.f (1/1)
beskattningenfinska (2/2)
därom (1/1)
arbetsliv (1/1)
förskoleenheter (1/1)
alakoulu (1/1)
sjukdagpenningfinska (2/2)
tänker (2/2)
fallit (3/3)
internetsidor (1/1)
vårdenhet (2/2)
företagstjänster (1/1)
kollektivavtalet (14/14)
församling (7/7)
klasserna (1/1)
identifieras (1/1)
konstuniversitet (2/2)
tidsbokningfinska (1/1)
grundskolanengelska (1/1)
brottmål (3/3)
frukter (1/1)
studieresor (1/1)
Bostadslöshet (1/1)
sakerna (1/1)
Mariegatan (1/1)
begravning (4/4)
familjehusen (1/1)
bokas (1/1)
båda (20/20)
utbildningssystemet (1/1)
österut (1/1)
ohälsa (1/1)
integritetsskydd (1/1)
närtågen (1/1)
ylletröja (1/1)
gynekologiska (2/2)
installera (1/1)
faderskapspenningdagar (4/4)
beviljande (1/1)
karneval (1/1)
lämpliga (2/2)
bekantar (1/1)
medling (6/6)
problemsituationer (1/1)
kvinnlig (2/2)
moderskapsförpackning (1/1)
polisstationen (6/6)
territorium (2/2)
finansieringsvederlag (1/1)
kompetensbaserat (2/2)
lov (1/1)
smidig (1/1)
fira (1/1)
frågar (2/2)
bevara (2/2)
grundare (2/2)
medborgarinstitut (8/8)
graviditetsintyg (1/1)
skuldrådgivningfinska (1/1)
elinkeinotoimisto (4/4)
företags (1/1)
företagarpensionsförsäkringenfinska (1/1)
chattenfinska (1/1)
hushållspapper (2/2)
arbetsplatsen (25/25)
handläggning (1/1)
hur (93/94) Hur (1)
absolut (1/1)
arbetsverksamhet (2/2)
korrekta (3/3)
ulkomaalaisten (1/1)
omfattande (6/6)
död (2/2)
utrikesministeriets (4/4)
placerar (2/2)
markägarens (1/1)
röster (2/2)
fots (2/2)
självrisken (2/2)
haku (1/1)
innevarande (1/1)
bostadsrättsbostadfinska (1/1)
Översättningar (1/1)
NTM (3/3)
lagstiftningen (6/6)
simhallar (4/4)
examensnivån (1/1)
erityishoitoraha (1/1)
säger (12/12)
Maahanmuuttajanuorten (1/1)
stödtjänster (6/6)
dialekterfinska (1/1)
Infobankens (3/3)
ensamstående (3/3)
ändrat (1/1)
volontärarbete (1/1)
konsulat (3/3)
lokaltrafikens (1/1)
ungdomsstationen (3/3)
tidtabeller (2/2)
lastensuojelu (1/1)
Lapset (1/1)
arbetsgivarförbunden (1/1)
anrika (1/1)
all (1/1)
yrkes- (2/2)
berör (5/5)
evenemang (9/9)
avlägga (56/56)
krisarbetare (1/1)
filmer (8/8)
fyllning (1/1)
förskoleundervisningenfinska (3/3)
bibehålla (2/2)
föreningsmedlemmar (1/1)
beredningen (1/1)
anmälningsblanketten (2/2)
frånvarande (2/2)
blankett (15/15)
snön (1/1)
graviditetsmånaden (5/5)
tidpunkt (2/2)
ansökningstiden (3/3)
utbildningfinska (2/2)
nyligen (5/5)
kansanopisto (2/2)
svenska (890/890)
ägda (1/1)
trygghet (13/13)
bostadsrättsbostäder (4/4)
studerandefinska (5/5)
resan (2/2)
tjänsteställe (11/11)
säljs (6/6)
besöket (3/3)
stjälande (1/1)
ordningsnummerfinska (1/1)
stödformer (1/1)
vigselhandlingarna (1/1)
samtalet (5/5)
bikulturellt (1/1)
äger (11/11)
skriftlig (7/7)
kommersiella (2/2)
förlovningen (1/1)
tjänsterfinska (9/9)
arbeten (1/1)
SIMHE (4/4)
begränsas (2/2)
mor- (4/4)
simma (1/1)
bemanningsbolag (1/1)
betonat (1/1)
suppleanter (1/1)
yttrandefrihet (1/1)
drabbats (1/1)
akademiska (1/1)
strax (1/1)
ombeds (1/1)
upphört (6/6)
ekonomiska (22/24) Ekonomiska (2)
publicera (1/1)
påsen (2/2)
YouTube (2/2)
springa (1/1)
högtidligt (1/1)
ägodelarna (1/1)
skiljas (3/3)
kräver (21/21)
undernivåer (1/1)
Österbotten (2/2)
hyresbostad (33/35) Hyresbostad (2)
personer (96/96)
farlig (1/1)
förvärvsarbetar (2/2)
ofrånkomliga (1/1)
namnändring (3/3)
förpackningen (1/1)
går (43/43)
referensramen (1/1)
biljettpriser (2/2)
förgiftats (1/1)
genast (9/9)
barnlöst (1/1)
nytta (5/5)
missbruksproblemfinska (2/2)
släkting (6/6)
dagvårdsavgifter (2/2)
kommun (19/19)
förvaltningsrätten (1/1)
berättigad (2/2)
badstränder (1/1)
svårare (4/4)
samhörighet (1/1)
inlärningsresultaten (1/1)
livsfara (2/2)
snabbare (3/3)
fortfarande (9/9)
öppnar (11/11)
Chydeniusfinska (1/1)
babyns (1/1)
föreningen (12/14) Föreningen (2)
felfri (1/1)
kontaktuppgifter (6/6)
brottet (1/1)
föreslå (2/2)
katastrofer (1/1)
tusen (2/2)
ålders- (1/1)
serviceställen (2/2)
sopsortering (1/1)
talet (15/15)
rumänska (12/12)
jourhavande (2/2)
heltidsstuderande (1/1)
undertrycka (1/1)
matematik (1/1)
Ammatilliseen (1/1)
föräldrarnas (10/10)
moderskapsunderstöd (6/6)
prövotid (1/1)
försvar (1/1)
fostran (18/21) Fostran (3)
exemplar (1/1)
planer (1/1)
folkpensionens (1/1)
uppstartsföretag (2/2)
klagar (1/1)
komplettera (2/2)
mån.-fre. (4/4)
tortyr (1/1)
regionförvaltningsverken (1/1)
skolelever (1/1)
arbetsintyg (12/14) Arbetsintyg (2)
mediciner (2/2)
populäraste (1/1)
botas (1/1)
databank (1/1)
länders (5/5)
Laureas (1/1)
villkoren (15/15)
familjeband (25/25)
jämlikhet (4/6) Jämlikhet (2)
överlåter (2/2)
pensionerna (3/3)
relativt (4/4)
ansökte (2/2)
pensionsärenden (1/1)
kvällen (4/4)
funderingar (1/1)
grammatikengelska (1/1)
lärandet (1/1)
diskrimineringen (1/1)
treårigt (2/2)
internationella (19/21) Internationella (2)
lättare (6/6)
hjälptelefon (3/3)
oikeusaputoimisto (4/4)
Kvinnokliniken (1/1)
verksamhetscenter (2/2)
varvid (1/1)
specialiserade (1/1)
vattenskada (5/5)
hårdaste (1/1)
tiden (25/25)
ansökningsförfarandena (1/1)
skolhälsovårdaren (4/4)
akademiskt (1/1)
ekonomiskt (4/5) Ekonomiskt (1)
badrum (1/1)
flyttat (9/9)
försöka (1/1)
livligare (1/1)
mobiltelefonens (1/1)
skötseln (6/6)
tågbiljetter (1/1)
invandrararbete (1/1)
Juristförbunds (2/2)
färdigt (2/2)
risker (2/2)
osuuskunta (1/1)
här (32/32)
vårdutgifterna (1/1)
vattenledningar (2/2)
arbetsprov (2/2)
försäkrad (3/3)
studerandehälsovården (2/2)
blödande (1/1)
hot (12/12)
ylioppilaskokeet (1/1)
Kaustby (2/2)
-kuntayhtymä (1/1)
nätbankkoder (1/1)
kielioppi (1/1)
Petikkos (1/1)
utrymme (1/1)
motioner (1/1)
tidigast (2/2)
ifrågavarande (4/4)
guldåldern (1/1)
efterlevande (2/2)
stödtjänsterna (2/2)
familjedagvårdare (7/7)
Lumon (2/2)
grundskolorna (1/1)
föras (2/2)
arbetarskyddsinspektioner (1/1)
moderskapsledigheten (5/5)
skatteprocent (6/6)
inbrottstjuvar (1/1)
så (63/63)
sjukförsäkringen (13/13)
hemmet (36/36)
visumansökningsblankett (1/1)
avgiftsfritt (3/3)
isländska (1/1)
familjeträning (1/1)
civil (2/2)
skyldig (10/10)
smärtlindring (1/1)
upplevelser (1/1)
flaggar (1/1)
funktionsnedsättning (7/7)
Trafiksäkerhetsverkets (1/1)
samråd (2/2)
semestrar (3/3)
januari (12/12)
framskrida (1/1)
avtalat (4/4)
återflyttarefinska (1/1)
hyreshusbolaget (1/1)
folks (1/1)
itsehoitolääke (1/1)
specialiserat (2/2)
seder (5/5)
godtagbara (1/1)
kulturella (1/1)
underskrift (2/2)
Hyresboende (1/1)
avgör (3/3)
hinner (3/3)
bistå (2/2)
bedöms (7/7)
brandsläckaren (1/1)
huvudstaden (2/2)
södra (5/5)
ry (16/16)
tingsrättfinska (2/2)
turism (4/4)
rådgivningspunkt (1/1)
kyrklig (2/2)
psykoterapeutens (1/1)
Foreigners (2/2)
födelse (10/10)
Gustav (3/3)
arbetarskyddsföreskrifterna (2/2)
godkänns (3/3)
pension (16/17) Pension (1)
vietnamesiska (7/7)
LUVA (3/3)
kejsaren (1/1)
religionsundervisningen (2/2)
traditionsarbetefinska (1/1)
Anonyymit (1/1)
avlägsnande (1/1)
förvaltningsmyndigheter (1/1)
Liechtenstein (12/12)
medborgarskapet (1/1)
familjeplaneringsrådgivningen (1/1)
tisdagar (3/3)
skattemyndigheten (3/3)
permanenta (2/2)
representera (1/1)
den (588/602) Den (14)
över (82/82)
Torggatan (1/1)
studieort (1/1)
brandvarnaren (2/2)
fysik (1/1)
vore (2/2)
förlossningen (18/18)
besvarar (2/2)
moderskapsledig (3/3)
inhämtat (1/1)
hälsovårdens (1/1)
självständighetsdagens (1/1)
förföljd (2/2)
hette (1/1)
tillståndsenheter (1/1)
utsätts (1/1)
Resultatenheten (1/1)
lösas (3/3)
identitetsbevis (8/8)
dyrast (1/1)
vandringfinska (1/1)
tillfrågas (1/1)
Oodi (2/2)
lö (1/1)
apteekki (1/1)
webblanketten (1/1)
förflyttningstillstånd (1/1)
livssituationen (1/1)
freden (1/1)
kuntoutussuunnitelma (1/1)
skala (1/1)
Sport (5/7) sport (2)
Jakobstad (2/2)
äta (1/1)
kullfallna (1/1)
äldre (14/19) Äldre (5)
yrkeshögskolorna (2/2)
efternamnen (1/1)
skidor (2/2)
underrättelse (2/2)
planeras (1/1)
socialskydd (1/1)
november (4/4)
tillgången (2/2)
hälsostationernas (2/2)
utvecklat (1/1)
ledighet (4/4)
varor (5/5)
centralsjukhuset (1/1)
Vionojafinska (1/1)
skogen (2/2)
hotar (9/9)
avlagt (38/38)
självrisktiden (2/2)
drogbruk (1/1)
arbetefinska (1/1)
krävs (32/32)
kriisipäivystys (3/3)
läroanstaltens (2/2)
Migrationsverketfinska (1/1)
nätbankskoder (4/4)
studentkårer (2/2)
Kyllönen (2/2)
förutsättningar (3/3)
integritetsskyddet (1/1)
humanitärt (1/1)
studiebyrå (1/1)
blanketter (1/1)
föregående (1/1)
stadslotsen (1/1)
stapelrättigheter (1/1)
kvadratmeter (2/2)
utbildningstiden (2/2)
låg (1/1)
flyktingens (1/1)
lapsikaappaus (1/1)
avloppet (1/1)
alltid (66/66)
vitas (1/1)
batteriinsamlingslådor (1/1)
Helsingin (5/5)
avsnitt (5/5)
säljer (9/9)
fisketillståndfinska (1/1)
nationalpark (2/2)
lokaltidningar (2/2)
nationernas (2/2)
Vardagslivet (1/1)
servicestyrcentral (1/1)
inflyttningen (2/2)
hälsotjänster (3/3)
avioliiton (2/2)
klienter (8/8)
inkomstrelaterade (5/5)
tolkar (2/2)
religiösa (10/10)
deltidsarbeta (1/1)
hösten (9/9)
minnas (2/2)
uppkommer (1/1)
barndomen (1/1)
arbetsavtalslagen (2/2)
inriktade (3/3)
skolgången (2/2)
företagarutbildning (4/4)
InfoFinland.fi (2/2)
tandläkarkontroll (2/2)
avvika (3/3)
administration (1/1)
krismottagningen (1/1)
servicenummer (1/1)
fingeravtryck (1/1)
föråldrade (1/1)
kompletteringsutbildning (1/1)
civilstånd (1/1)
månadsskift (1/1)
jämföra (4/4)
vårdfinska (1/1)
rörelsehandikappad (1/1)
sjukhusen (1/1)
regel (7/7)
gången (2/2)
regelbundna (3/3)
lämnats (3/3)
samlat (1/1)
frivilliga (4/4)
fritidsaktiviteterna (1/1)
läkarremiss (2/2)
konsumentens (3/3)
hälsovårdsministeriet (3/3)
mellanmål (1/1)
kulturhistorisk (1/1)
ordnar (66/66)
företedde (1/1)
psykiatrian (1/1)
ansluta (10/10)
idrottsplaner (2/2)
invandrare (86/86)
perhehoito (1/1)
avbokar (1/1)
högsommarens (1/1)
enheten (4/4)
kommunalskatt (1/1)
faderskap (4/4)
torsdag (2/2)
lampor (2/2)
säga (23/23)
bibliotekstjänstfinska (1/1)
alternativ (8/8)
snart (1/1)
tryggat (2/2)
tjänsterna (31/31)
undervisningfinska (2/2)
sköta (21/21)
trivas (1/1)
kotivakuutus (1/1)
verksamhetsformerna (1/1)
tryggheten (61/61)
följaktligen (1/1)
Konsumentrådgivningen (1/2) konsumentrådgivningen (1)
borgerliga (1/1)
språkcaféerna (2/2)
ni (42/42)
tjänsten (64/64)
lyhytkurssi (1/1)
skrivs (4/4)
utfärdad (1/1)
civiltjänstgörare (2/2)
tidpunkten (5/5)
hemvårdsstödet (3/3)
beaktar (2/2)
sjukvårdskostnader (2/2)
ålderdom (1/1)
arbetsgivarförbundet (1/1)
nationalspråk (2/2)
konflikterna (2/2)
bostadssidor (1/1)
kommunikation (4/4)
månatliga (1/1)
uppehållsrätten (18/18)
hyrt (1/1)
bibliotek (16/17) Bibliotek (1)
gymnasieskolor (2/2)
blanketten (18/18)
möjligheter (11/11)
bostadslån (7/7)
ärendena (1/1)
bostadsaktiebolag (5/5)
mäklararvode (1/1)
nästan (12/12)
vanligt (9/9)
mål (3/3)
sammanträden (3/3)
stöder (8/8)
väst (2/2)
hissa (1/1)
Karlebyfinska (5/5)
psykiskt (1/1)
inverkar (6/6)
dagpenningen (4/4)
industrialiserades (1/1)
belopp (23/23)
förtroendeuppdrag (1/1)
hårt (1/1)
mörkt (1/1)
Vasa (6/6)
kartläggningfinska (1/1)
invid (1/1)
omavastuuaika (2/2)
InfoFinland (21/21)
förmånligast (1/1)
kreditgivning (1/1)
tillståndsärenden (4/4)
originalhandlingen (1/1)
webbapotek (1/1)
ange (8/8)
fortsättningsvis (1/1)
förlorat (1/1)
bokbussar (1/1)
tag (1/1)
skapa (7/7)
käräjäoikeus (3/3)
Karl (1/1)
president (4/4)
sörja (4/4)
mamma- (1/1)
Finnvera (3/3)
sorani (3/3)
texttelefon (1/1)
förnyas (1/1)
webbtjänster (2/2)
banker (3/3)
betraktats (1/1)
även (347/347)
infödd (4/4)
höra (5/5)
problemfinska (2/2)
studiestödetengelska (1/1)
asunnot (6/12) Asunnot (6)
åldersgränser (1/1)
missbruk (2/2)
trafikförsäkring (1/1)
tillkalla (1/1)
fördel (2/2)
pepparkakor (1/1)
Migrationsverkets (27/27)
inhemska (3/3)
rimliga (1/1)
studerat (3/3)
förmåner (28/28)
råd (89/89)
affären (1/1)
OYS (1/1)
ersättas (1/1)
Akava (1/2) AKAVA (1)
textade (1/1)
lokaltidningen (3/3)
särskild (6/6)
hittar (202/202)
undervisar (4/4)
penningunderstödfinska (1/1)
kortare (5/5)
medlem (20/20)
medborgarskap (70/70)
levt (1/1)
familjepensionsskydd (1/1)
badrumsrenovering (1/1)
synskadadefinska (1/1)
verksamhetsplanen (1/1)
upphörande (2/2)
prioriteten (1/1)
beskattningsbeslutfinska (1/1)
Kehitysvammaliittos (1/1)
jämte (1/1)
Gammelstadsforsen (1/1)
identifiering (2/2)
övervakar (10/10)
sammanställts (1/1)
Studenternas (1/1)
centralerna (1/1)
snabel (1/1)
straffpåföljd (1/1)
internationellt (8/8)
medelhög (1/1)
skattepengar (1/1)
diskriminerings- (2/2)
Advisor (1/1)
sjukhusvård (2/2)
yngsta (2/2)
samhällsvetenskapliga (3/3)
med (667/667)
skolors (1/1)
följeslagare (1/1)
inkomster (34/34)
förbinder (1/1)
förpackningsmaterial (1/1)
tandvårdstjänster (1/1)
källskatt (1/1)
kyrkoherden (1/1)
specialyrkesläroanstalter (1/1)
SHVS (1/1)
boendefrågor (1/1)
garantin (1/1)
spanska (37/37)
seudun (3/3)
årskurser (1/1)
barnpassningsservicen (1/1)
atmosfär (1/1)
Vandakanalen (1/1)
bostadsrätten (2/2)
beskickning (16/16)
folkmängd (1/1)
temperaturerna (1/1)
hemkommuns (3/3)
används (7/7)
branschen (2/2)
U2 (1/1)
pågå (1/1)
hälften (1/1)
poliklinik (1/1)
fadern (10/10)
simhallen (1/1)
dagvårdsplatser (1/1)
medelst (2/2)
brottsanmälan (7/7)
anknutna (1/1)
jobbansökan (5/5)
begå (2/2)
rådgivning (54/54)
användande (1/1)
passfoto (2/2)
ansökningar (4/4)
välgrundad (3/3)
handelsstad (2/2)
åldrar (5/5)
väljas (4/4)
fastighetsförmedlare (1/1)
koppling (1/1)
gifter (4/4)
Matkahuoltos (4/4)
specialyrkesexamen (3/3)
teckenspråkstolk (1/1)
uppge (5/5)
stadshuset (2/2)
laga (3/3)
kyrkans (3/4) Kyrkans (1)
tull- (1/1)
återvinns (1/1)
åldringar (4/4)
studiebetyg (1/1)
ändringsarbeten (2/2)
specialvårdpenning (2/2)
ingenjör (1/1)
blåser (1/1)
tillhandahåller (19/19)
handlägger (1/1)
konsumenter (1/1)
växande (1/1)
studievägledarna (2/2)
begravningsplatser (4/4)
hårdare (1/1)
efterhand (5/5)
utfärder (2/2)
motiverade (1/1)
nättjänst (1/1)
införde (2/2)
upplevs (1/1)
intervjuar (1/1)
registrera (36/36)
Lichtenstein (1/1)
skogsbruksområden (1/1)
långtidssjuka (2/2)
föräldern (23/23)
mark (3/3)
fruktar (2/2)
kommunvalfinska (1/1)
befolkning (2/2)
viken (3/3)
central (2/2)
temperaturen (2/2)
låna (10/10)
välbefinnande (1/1)
näringstjänsterfinska (2/2)
förskoleplats (4/4)
ansökningssättet (1/1)
webbsidan (1/1)
ansvar (8/8)
kursavgiften (2/2)
RAMK (2/2)
dagvården (13/13)
rehabiliteringspenning (2/2)
nybörjarkurser (1/1)
lisä (1/1)
rusmedelsmottagning (1/1)
marknadsundersökning (1/1)
kan (1874/1875) Kan (1)
fastställts (5/5)
följeslagartjänstfinska (2/2)
Marthaförbundet (1/1)
materialet (4/4)
riksdagenfinska (1/1)
V (2/2)
läsårsavgiften (2/2)
företagsformerfinska (1/1)
hembygdsmuseer (1/1)
uppringd (2/2)
medicinsk (13/13)
deltidsarbete (1/1)
därefter (12/12)
vokabulär (2/2)
förpackningar (3/3)
medlare (2/2)
jokamiehen (1/1)
familjerna (1/1)
socialväsen (2/2)
utlandetfinska (1/1)
frånvaro (1/1)
studiemiljö (2/2)
nödcentralen (2/2)
affärsverksamhet (3/3)
startpaket (1/1)
kö (1/1)
lönsam (3/3)
sidoapotek (1/1)
Kafnettis (1/1)
Ylikylä (1/1)
perustamisilmoitus (1/1)
på (1686/1687) På (1)
värmesystem (1/1)
Nordisk (3/4) nordisk (1)
blir (59/59)
förskolan (4/4)
straffas (1/1)
elev- (1/1)
alle (1/1)
elavtal (4/4)
öarna (2/2)
välbefinnandeområden (1/1)
hallen (1/1)
arbetstiderna (1/1)
Mellersta (11/13) mellersta (2)
be (44/44)
hälsovårdstjänsterna (21/21)
papperslöshetfinska (1/1)
borgen (6/6)
fyrverkerierna (1/1)
fördelas (1/1)
kursernas (1/1)
inskrivet (1/1)
läroanstalter (17/17)
läroavtalsbyrån (1/1)
lindras (1/1)
gruppen (5/5)
familjen (49/49)
dagvårdsplatsfinska (2/2)
flygresor (1/1)
vigselintyg (1/1)
omfattning (5/5)
verksamma (5/5)
utanför (17/17)
premier (1/1)
kunden (6/6)
flickorfinska (2/2)
väst- (2/2)
börjar (34/34)
rättegång (1/1)
Musikantitfinska (1/1)
humanistiska (4/6) Humanistiska (2)
mall (1/1)
redan (30/30)
inkomsten (2/2)
entreprenörskap (5/5)
abikurssi (1/1)
annonserar (1/1)
pengarna (1/1)
fiskelov (1/1)
säljaren (7/7)
Opetushallitus (5/7) opetushallitus (2)
ennakonpidätys (2/2)
bönestund (1/1)
samtal (4/4)
Garantistiftelsen (1/1)
semesterresa (1/1)
mötesplatsen (1/1)
vuotiaan (1/1)
högersinnade (1/1)
upprätthållande (1/1)
ansökningsproceduren (1/1)
begränsningarna (4/4)
skor (1/1)
självständig (2/2)
köket (1/1)
ungdomsfullmäktige (1/1)
informering (1/1)
bostadslös (3/3)
bibliotekarien (2/2)
krävas (1/1)
lärt (3/3)
ej (1/1)
psykiatriska (1/1)
blivit (30/30)
avslå (1/1)
tillhörande (1/1)
kommunfinska (1/1)
nödcentraloperatörens (1/1)
betalades (2/2)
välhållen (1/1)
Karlebynejdens (2/2)
sairaala (2/2)
valuta (4/4)
vaarallinen (1/1)
naturstigar (1/1)
vuxen (5/5)
offentliga (56/56)
koordinatoren (1/1)
utkomstskyddet (4/4)
F (1/1)
dammsugaren (1/1)
narkomaner (2/2)
allmänbildande (3/3)
kollegor (3/3)
autovero (1/1)
någondera (3/3)
landskapsmuseumfinska (1/1)
daggymnasiet (1/1)
fotot (1/1)
utfärdats (10/10)
prövas (2/2)
sedan (11/11)
vetenskaplig (1/1)
elektriska (2/2)
offer (24/24)
arbetstagaren (16/16)
samtalsklubbar (1/1)
verkets (1/1)
ofta (44/44)
minimivillkor (1/1)
informerar (5/5)
vilket (44/44)
hon (47/47)
uträtta (3/3)
kalla (2/2)
landsvägsförbindelsermed (1/1)
vite (1/1)
fristående (9/9)
högteknologiska (1/1)
hyresbostäderengelska (1/1)
kandiderar (1/1)
fastighetsskötseln (3/3)
moderskapspenning (9/9)
ringer (13/13)
programmet (1/1)
Romppu (1/1)
färdmedel (1/1)
gäller (40/40)
intresse (4/4)
evenemangskalenderfinska (1/1)
Internetanslutningar (1/1)
Rovaniemi (42/42)
överenskommelsen (3/3)
Handelsbanken (1/1)
Infobanken (5/5)
bryter (4/4)
yrkeshögskoleexamen (10/10)
summa (4/4)
Tavastehus (1/1)
automatik (1/1)
filmerfinska (1/1)
kotihoidon (2/2)
finsk- (1/1)
hälsovården (18/18)
d.v.s. (14/14)
paddling (1/1)
böckerna (1/1)
drag (1/1)
historiafinska (1/1)
mottagit (1/1)
kontakta (116/116)
Kaapatut (1/1)
fördelningen (3/3)
Helsingforsregionen (5/5)
bokföringen (6/6)
gravkvarter (1/1)
perustoimeentulotuki (1/1)
uppskattning (2/2)
ersättningsgilla (1/1)
nämna (1/1)
produkt (1/1)
flicka (1/1)
Kompetenscentret (1/1)
matka.fi (1/1)
uppehållstillstånd (269/274) Uppehållstillstånd (5)
utbildningskoncernfinska (1/1)
såvida (1/1)
rum (4/4)
minnesproblemen (1/1)
informations- (2/2)
hembesök (2/2)
områdeskoordinatorn (1/1)
tåg- (1/1)
skyddshuset (1/1)
antagen (4/4)
hälsorådgivningen (2/2)
elatustuki (1/1)
korrigerar (1/1)
universitetsutbildningfinska (1/1)
vardagsmotion (1/1)
Räckhals (1/1)
resedokumentfinska (1/1)
fortsatt (13/15) Fortsatt (2)
webbaserade (1/1)
utbetalat (1/1)
föräldradagpenningens (1/1)
Fpas (1/1)
maskinmästare (1/1)
kunde (2/2)
änka (2/2)
avstängda (1/1)
utexaminerats (1/1)
esiopetus (3/3)
kläder (6/6)
oleskelulupa (1/1)
minns (4/4)
kunderna (10/10)
självrisktid (2/2)
bostadsrättsavtalet (1/1)
hälsorisk (1/1)
parförhållanden (3/3)
utgångsläge (1/1)
tid (148/148)
Nylands (10/10)
läsning (2/2)
hålls (8/8)
annan (65/65)
asylprocessens (1/1)
möte (5/5)
medför (1/1)
församlings (3/3)
godta (1/1)
Helsingforsregionen.fi (1/2) HelsingforsRegionen.fi (1)
uppfattning (1/1)
boendet (9/9)
extra (4/4)
tull (1/1)
MinSkatt (3/3)
civiltjänstgöring (1/1)
vuxenutbildningsinstitut (4/4)
ingripa (3/3)
måltidsstödet (1/1)
inträdesprov (2/2)
dygnet (25/25)
skridskobanor (1/1)
bostäderfinska (2/2)
servicerådgivning (1/1)
Peijaksen (2/2)
Kiasmafinska (1/1)
nationalparker (1/1)
servicehandledning (1/1)
semesterna (1/1)
bärande (1/1)
tar (52/52)
tätskikt (1/1)
sjukhuskostnaderna (1/1)
betalas (44/44)
Spafinska (2/2)
äktenskapengelska (1/1)
installeras (1/1)
samtidigt (25/25)
Huvudstadens (3/3)
länken (3/3)
idkar (1/1)
bedrivs (1/1)
lämnade (4/4)
garanti (2/2)
sysselsättnings- (1/1)
slag (2/2)
bosättning (2/2)
före (52/52)
utbildningar (7/7)
tidsbestämt (8/8)
värdefull (1/1)
bett (2/2)
palvelutalo (1/1)
utkommer (3/3)
säsongsarbete (2/2)
möjligheten (3/3)
neuvola (4/4)
arbetstillstånd (1/1)
ålderspension (5/5)
polska (13/13)
livsmiljö (1/1)
söker (41/41)
ehkäisyneuvola (1/1)
slut (4/4)
förbereda (2/2)
framtid (2/2)
säkerställa (5/5)
avstånd (1/1)
markägaren (1/1)
onyktert (1/1)
konflikter (5/5)
fortsatte (1/1)
partiell (9/9)
sin (75/75)
kontrakt (1/1)
handikappbidrag (5/5)
redogörelsen (1/1)
kontot (1/1)
ositus (1/1)
förskrivningsrätt (1/1)
arbetarinstitutets (1/1)
stiger (4/4)
klarlägga (1/1)
videkvistar (1/1)
kompletteras (2/2)
midsommar (1/1)
säkerhet (11/11)
näringsidkande (1/1)
kunskapscenter (1/1)
grannländer (2/2)
kosta (1/1)
elev (2/2)
kortfattade (1/1)
lekverksamhet (1/1)
FöretagsEsbo (1/1)
Skatteförvaltningen (4/5) skatteförvaltningen (1)
föräldrarna (51/51)
krissituation (5/5)
lyckades (2/2)
baserat (4/4)
yhteispäivystys (1/1)
ordböckerfinska (2/2)
kulturförening (1/1)
bearbetningar (1/1)
bilder (3/3)
förhöjningsdelen (1/1)
flertal (1/1)
barnrådgivning (1/1)
medeltalet (1/1)
Internetuppkoppling (1/1)
krishjälp (1/1)
maximibelopp (1/1)
läkarintyg (5/5)
handledningstjänster (1/1)
invånarantal (1/1)
caféer (1/1)
kommunaval (1/1)
kundtjänst (1/1)
lång (17/17)
höga (1/1)
pålitligt (3/3)
djuren (1/1)
massörexamen (1/1)
befolkningsdatasystemet (14/14)
hjälptelefonen (2/2)
stadigvarande (45/45)
skjuta (1/1)
tillåtna (2/2)
oikeusturvavakuutus (1/1)
linkkiFörsamlingen (1/1)
verkosto (1/1)
invånarverksamheten (1/1)
bestämda (1/1)
perukirja (1/1)
Akatemia (3/3)
bildkonstskola (1/1)
ersättningen (1/1)
vänta (8/8)
hörselnfinska (1/1)
kaffe (1/1)
Haag (1/1)
vuokrasopimus (1/1)
godkännas (1/1)
Barnskyddsförbund (4/5) barnskyddsförbund (1)
utbildningsprogram (8/8)
utvecklingsstördafinska (1/1)
branscher (10/10)
det (475/476) Det (1)
enfas (2/2)
mödrar (1/1)
sommarsolståndet (1/1)
Eiran (1/1)
ovan (4/4)
konto (13/13)
hörselundersökning (1/1)
familjemedlemmar (21/21)
förskottsskatt (1/1)
huvudstadsregionen (12/12)
aktiveringsmodellen (1/1)
part (5/5)
utförs (4/4)
står (11/11)
studentbostadsstiftelse (6/6)
syften (1/1)
samhällsmedlem (1/1)
intresseorganisationfinska (1/1)
dessafinska (1/1)
drogproblemfinska (1/1)
jourtelefonen (2/2)
samfund (17/17)
klockslaget (1/1)
advokat (1/1)
halvvägs (1/1)
Salutorget (1/1)
taxa (1/1)
samhällelig (1/1)
högre (26/26)
gårdsområdet (1/1)
tidsperioder (1/1)
nuorisopsykiatrian (1/1)
uppgår (1/1)
inlärningssvårigheter (1/1)
begränsad (4/4)
hälsafinska (2/2)
kvarter (1/1)
marknadsföring (1/1)
tvisten (1/1)
byggplats (1/1)
påse (1/1)
gärna (3/3)
lunchsedlar (1/1)
officiellt (11/15) Officiellt (4)
universitetet (19/19)
intyget (11/11)
mottagningscenter (1/1)
arbetserfarenheten (1/1)
grundas (3/3)
diskrimineringfinska (1/1)
delägarbostad (2/3) Delägarbostad (1)
ingå (10/10)
förflutit (1/1)
bokar (11/11)
hotfull (1/1)
kierrätys.info (1/1)
utförandet (5/5)
gymnasiumfinska (1/1)
förverkligas (3/3)
munhälsovårdfinska (1/1)
lyftanordningar (1/1)
taitavan (1/1)
Finland (1008/1008)
perioden (2/2)
närstående (20/20)
biogas (1/1)
privatpersoners (1/1)
Simundervisnings- (1/1)
släkten (1/1)
hälsostations (1/1)
familjerådgivningsbyråerna (1/1)
söndagen (1/1)
folkpension (6/6)
Kafnetin (1/1)
följande (48/48)
fattas (10/10)
väljs (12/12)
uppstartsföretagare (11/11)
fortsätta (8/8)
livmodern (1/1)
utkomst (6/6)
Håkansböle (6/6)
enkel- (1/1)
underhålls (1/1)
uppfattas (1/1)
val (13/16) Val (3)
vårdande (1/1)
tvåspråkiga (4/4)
teknisk (1/1)
MoniNets (4/4)
oåterkalleligt (1/1)
näringslivstjänsterna (1/1)
in (81/85) In (4)
populärare (1/1)
adress (27/27)
livskompetensen (1/1)
grundval (1/1)
förhållandet (1/1)
hemlig (1/1)
väntat (1/1)
smarttelefonen (1/1)
moderskapspenningperioden (1/1)
faktum (1/1)
förläggning (1/1)
Klockarmalmens (1/1)
lisensiaatti (1/1)
tapaturmavakuutus (1/1)
arbetsamhet (1/1)
bortföranden (1/1)
historiska (4/4)
lastenvalvoja (3/3)
obligatorisk (2/2)
turism- (2/2)
sysslor (1/1)
rehabiliteringar (1/1)
lågstadiet (2/2)
stadgade (1/1)
kejsare (1/1)
studiepenningens (1/1)
växelverkan (2/2)
VALMA (13/13)
hemförsäkring (5/5)
födelsen (1/1)
museot.fi (1/1)
umgänge (2/2)
bikulturella (1/1)
lek (2/2)
företagarutbildningar (1/1)
kommersiellt (1/1)
genomsnittliga (1/1)
passfinska (1/1)
språkkaféer (1/1)
peruspäiväraha (1/1)
allvarlig (1/1)
kulturer (6/6)
avfallshanteringen (1/1)
tillgänglig (2/2)
enligt (53/53)
gymnasiestudierfinska (1/1)
uppmuntras (1/1)
ingreppet (1/1)
förkortat (1/1)
varsel (1/1)
underhållsskyldigafinska (1/1)
tydlig (1/1)
e (29/30) E (1)
nordligaste (2/2)
skuldlinjen (1/1)
personförsäkring (1/1)
hyresbostäder (32/32)
arbetstagarna (3/3)
hobbyverksamheter (2/2)
brottsmål (1/1)
resa (7/7)
förorsakat (1/1)
brand (9/9)
syfte (2/2)
herraväldet (1/1)
luthersk (1/1)
äter (4/4)
köpeanbudet (2/2)
tillbaka (6/6)
tukipiste (2/2)
beslutsfattandet (6/6)
byråerfinska (1/1)
vuxengymnasium (12/13) Vuxengymnasium (1)
gemensamt (11/11)
skattefritt (1/1)
inkomstrelaterat (1/1)
Ungdomspolikliniken (1/1)
sommar- (1/1)
försörjer (1/1)
förmiddagar (1/1)
holländska (10/10)
fyll (4/4)
separeras (1/1)
närserviceprincipen (2/2)
HelsingforsHels (1/1)
påverkar (14/14)
utrymmen (1/1)
funktionsförmågan (2/2)
hamnat (2/2)
lekar (1/1)
ansökningsblanketten (3/3)
idrott (3/3)
filmvisningarfinska (1/1)
penningspelproblemfinska (1/1)
tagalog (1/1)
läser (8/8)
rör (40/40)
konkurrera (1/1)
hygienföreskrifter (1/1)
sjukskrivning (1/1)
Spektr (1/1)
skötsel (2/2)
uttryck (2/2)
arbeta (80/82) Arbeta (2)
läroanstalt (12/12)
fulla (1/1)
Folkmusik (1/1)
många (143/143)
Setlementti (7/7)
Valviras (1/1)
pensionssystemen (1/1)
tema (1/1)
verkligen (3/3)
reseplanerare (1/1)
bilteknik (1/1)
öva (2/2)
gångfinska (1/1)
fås (14/14)
verifiera (1/1)
löfte (1/1)
lagarfinska (1/1)
utgång (1/1)
sägs (1/1)
vården (11/11)
yrkesläroanstalt (8/8)
ansvarsområde (1/1)
flykting (8/9) Flykting (1)
Ruokavirasto (1/1)
hemlands (4/4)
chefredaktör (2/2)
låta (7/7)
om (1845/1851) Om (6)
besökare (1/1)
Folkdans (1/1)
finskakurs (1/1)
camping (1/1)
Dickursby (4/4)
kollektivavtal (4/4)
Nyföretagarcentral (1/1)
idrottsklubbar (6/6)
PUK (1/1)
stora (15/16) Stora (1)
portugisiska (18/18)
renkött (1/1)
eftermiddagen (2/2)
ärendet (11/11)
avsikt (2/2)
språketengelska (1/1)
museikvarterens (1/1)
värdesätter (3/3)
hätänumero (2/2)
filmens (1/1)
kvällar (6/6)
gränsen (1/1)
stickkontakt (1/1)
Ristrand (1/1)
problemet (1/1)
misstag (1/1)
förfaringssätten (1/1)
könssjukdom (3/3)
rådgivningstelefon (1/1)
meningar (1/1)
bidragen (1/1)
boendekostnader (5/5)
betalningssvårigheter (1/1)
personuppgifter (5/5)
utredning (15/15)
dras (4/4)
AA (2/2)
hela (27/27)
Suomessa (2/2)
anhöriga (10/10)
bok (1/1)
löften (1/1)
karensen (1/1)
vardagliga (4/4)
vårdsystemet (1/1)
ha (119/119)
brottfinska (1/1)
medborgarorganisationer (1/1)
bodelningen (4/4)
integrationsutbildning (5/5)
välfärd (6/6)
upptäcker (8/8)
aktörerna (1/1)
konkreta (1/1)
ammattiopisto (4/4)
daghem (34/34)
oroar (1/1)
ogiltigt (1/1)
sjukvården (11/11)
tillstånd (57/57)
sysselsättningen (1/1)
InfoFinlands (289/289)
polisen (18/19) Polisen (1)
skolresor (1/1)
personlig (8/8)
dateras (1/1)
lönearbete (3/3)
fastställa (1/1)
dubbelnamn (1/1)
återförenas (1/1)
dyrare (11/11)
grundlagenfinska (1/1)
medverkar (2/2)
midsommareldar (1/1)
asylansökanfinska (1/1)
EU:s (2/2)
vilken (39/39)
sexuella (6/6)
förmodligen (1/1)
rubrik (1/1)
byggnaderna (1/1)
jag (54/54)
asyl (20/20)
ehkäisy (1/1)
regiontaxi (1/1)
bostadsbehov (4/4)
flygstationen (1/1)
önskemål (6/6)
utlänning (2/2)
tryggare (1/1)
intressebevakning (1/1)
familjerådgivningen (18/18)
sjukförsäkringsersättningen (1/1)
Avfallshantering (3/4) avfallshantering (1)
inslag.Om (1/1)
barnlöshet (1/1)
Helsinki (11/11)
född (1/1)
tidtabellen (1/1)
arbetsförhållanden (3/3)
bero (1/1)
tjänstekollektivavtalet (1/1)
kvinnans (2/2)
sätta (1/1)
utlämnad (1/1)
examensinriktad (1/1)
sosiaali- (4/6) Sosiaali- (2)
lös (1/1)
enskild (4/4)
fastställt (1/1)
Sato (2/2)
funktionalitet (1/1)
småbarnsfostran (4/4)
arbetslagstiftningen (2/2)
semesterpenning (1/1)
Tullen (1/1)
lånord (1/1)
restaurang (3/3)
diabetes (2/2)
möjliga (1/1)
enheter (2/2)
behålla (1/1)
betalat (10/10)
ersättningar (1/1)
sommartid (1/1)
sidor (18/18)
studietid (1/1)
juristens (1/1)
30l (1/1)
färre (1/1)
Chydenius (2/2)
velkaneuvonta (1/1)
kulturhus (1/1)
äe (1/1)
vattenkranarna (1/1)
Kronoby (1/1)
Monika (3/3)
betalda (1/1)
biografkedjan (1/1)
eleverna (5/5)
studielivet (1/1)
klarar (11/11)
gymnasierna (2/2)
arbetar (40/40)
fredag (8/8)
japanska (6/6)
allmännyttiga (1/1)
sjukpenning (1/1)
varje (35/35)
länderna (18/18)
publikationer (1/1)
övertid (2/2)
länk (3/3)
cookies (1/1)
exporterade (2/2)
mig (3/3)
rättelserna (2/2)
linkkiLaNuti (1/1)
makten (4/4)
boenderådgivare (1/1)
familjeledigheten (2/2)
samarbetsavtal (2/2)
söka (138/138)
kväll (1/1)
rätta (4/4)
motionsform (1/1)
centralsjukhus (3/3)
Sanomat (1/1)
arbetserfarenhet (10/10)
bollplaner (1/1)
yrkeshögskoleexamina (1/1)
förbundet (2/3) Förbundet (1)
skolgångsbiträde (1/1)
invandrartjänster (1/1)
nyfödda (1/1)
utrikes (1/1)
jobbsajterfinska (1/1)
sjukdagpenningen (3/3)
sökordet (1/1)
välkomna (3/3)
behovsprövad (3/3)
beskattningsrätt (1/1)
affärer (1/1)
människohandelns (2/2)
ledigheterna (1/1)
negativt (4/5) Negativt (1)
fullt (1/1)
pilkning (1/1)
lähetetty (1/1)
eleven (2/2)
Reittiopas (2/2)
Rovalan (7/7)
överenskommelse (3/3)
förrätta (1/1)
Centria (1/1)
stort (8/8)
rehabiliterande (2/2)
läroanstalternas (2/2)
katolska (2/2)
bostäderna (4/4)
samarbete (4/4)
väljer (10/10)
fadernfinska (1/1)
kontaktspråket (1/1)
vistelsen (4/4)
traditioner (1/1)
arkitektur (2/2)
meddelas (8/8)
tingsrätt (3/3)
påbrå (1/1)
maistraatti.fi (2/2)
miljon (1/1)
grundlagfinska (1/1)
skol- (1/1)
snö (1/1)
kommande (1/1)
knappsatsen (1/1)
utlänningars (1/1)
ansvaret (9/9)
arbetarinstituten (2/2)
inkassobyrån (1/1)
arbetsgivare (63/63)
kommuntillägg (4/4)
höger (1/1)
KOSEKs (1/1)
syrjintä (1/1)
ordentlig (2/2)
baseras (1/1)
Livräddningsförbund (1/1)
våldsamt (3/3)
ikäihmisten (1/1)
djur (1/1)
Mielenterveysseura (3/3)
uppdragsgivare (1/1)
lyckas (1/1)
antagningen (1/1)
slås (1/1)
behövs (28/28)
svenskan (2/2)
slidmynning (1/1)
förtjänade (1/1)
Ounasälv (1/1)
utbildningen (53/53)
registreras (20/20)
internetionellt (1/1)
visumfritt (2/2)
fått (44/44)
säkerheten (3/3)
vårdnadshavarens (1/1)
turneringar (1/1)
läkemedelsförpackningen (1/1)
införskaffat (1/1)
främmande (9/9)
hurdant (4/4)
beloppet (5/5)
reservera (4/4)
inkomstgräns (1/1)
palveluasuminen (1/1)
tvätt- (1/1)
mekanisk (1/1)
detta (95/95)
rösträttsregistret (6/6)
medlemsland (1/1)
vän (7/7)
kombinerat (5/5)
yhdenvertaisuus (1/1)
Iso (5/5)
försäkringsintyg (1/1)
postfack (1/1)
stipendier (4/4)
lider (2/2)
eld (2/2)
bereder (2/2)
dröjsmål (1/1)
asukastila (1/1)
snöar (1/1)
efteråt (1/1)
flexibel (7/7)
kund (12/12)
familjeledighet (2/4) Familjeledighet (2)
koululaisten (1/1)
vederlag (2/2)
slottets (1/1)
Lumo (1/1)
kiosker (4/4)
bär (4/4)
nu (1/1)
hade (7/7)
Schengenvisumfinska (1/1)
fruktan (1/1)
kulturministeriet (4/4)
trafikreglerna (2/2)
självfinska (2/2)
närmare (13/13)
logi (1/1)
utfärdar (2/2)
format (4/4)
estetiska (1/1)
självständigt (14/14)
HRT (3/3)
ungefär (16/16)
lokaltrafik (1/1)
bibliotekskort (7/7)
webbsidorna (1/1)
läroplikt (3/3)
Turku (1/1)
starttiraha (1/1)
handikappat (8/8)
undersökas (1/1)
sammanfattning (3/3)
magistraten (87/88) Magistraten (1)
stadgarna (1/1)
Inkomstregistret (1/1)
utbetalningen (2/2)
underuthyrning (1/1)
delaktig (1/1)
förman (1/1)
morgon (2/2)
webbplatsen (19/19)
Sveaborg (2/2)
utarbeta (3/3)
tillståndsärende (1/1)
plastförpackningarna (1/1)
invandrares (2/2)
Alberga (1/1)
arbetarinstitut (11/11)
översättning (1/1)
tilläggsundervisning (2/2)
frånskild (1/1)
dagvårdstjänster (2/2)
ugnen (1/1)
tionde (5/5)
svårigheter (3/3)
idrottsanläggningar (1/1)
förändras (1/1)
Seniorinfo (1/1)
servicerådgivare (1/1)
tjära (3/3)
lokalförvaltningfinska (1/1)
trafikknutpunkt (1/1)
styr (1/1)
redaktör (1/1)
huruvida (7/7)
översättare (4/4)
ansökning (5/5)
för (1620/1622) För (2)
gren (1/1)
arbetslöshetskassa (9/10) Arbetslöshetskassa (1)
letar (5/5)
arbetspensionsanstalten (3/3)
mobiltelefontillverkaren (1/1)
bisyssla (2/2)
officiella (5/5)
norska (9/9)
byggd (1/1)
grupper (11/11)
yrkeshögskolafinska (3/3)
P (3/5) p (2)
vardagsum (1/1)
utarbetandet (1/1)
regelbunden (2/2)
tyst (3/3)
engelskspråkiga (3/3)
Dövas (3/3)
nutidskonst (1/1)
städa (1/1)
Kivenkolo (5/5)
Grani (2/2)
paret (2/2)
ekonomin (1/1)
god (11/12) God (1)
behandling (9/9)
felen (1/1)
viktigt (30/30)
Infobank (1/1)
doseras (1/1)
anställningsförhållande (1/1)
områdets (2/2)
faderskapsledighet (3/3)
belagt (1/1)
människor (37/37)
ju (1/1)
konsthusen (1/1)
telefontjänsten (6/6)
offret (1/1)
rekreationsdagar (1/1)
arbetarskyddschef (1/1)
applikationer (1/1)
Kokkolan (1/1)
ASE (7/7)
bibliotekfinska (1/1)
Lapplands (21/21)
ungdomsväsende (1/1)
tillgängligheten (1/1)
myndigheterfinska (1/1)
Österbottens (17/17)
for (2/2)
kontinuerliga (3/3)
överallt (1/1)
demonstrationer (1/1)
flyktingen (1/1)
webbtjänstfinska (1/1)
religionsutövande (1/1)
finansierade (3/3)
betänketid (2/2)
intresserad (8/8)
hyresgästen (4/4)
något (71/71)
adoptera (1/1)
dött (2/2)
joggingbanor (1/1)
hemhjälpfinska (1/1)
läsa (16/16)
säljas (1/1)
partnern (2/2)
eKirjasto (1/1)
östra (2/3) Östra (1)
skötandet (2/2)
socialbyrå (2/2)
familjerådgivningfinska (1/1)
enhet (7/7)
typer (4/4)
medlas (1/1)
assistentens (1/1)
Celsiusgrader (3/3)
Infopankki.fi (1/1)
yhdenvertaisuus- (1/1)
elledningar (2/2)
flyktingbakgrund (1/1)
&quot; (14/14)
preventivmetoder (1/1)
graviditetenfinska (1/1)
närmaste (20/20)
tillvalsämnen (1/1)
jämkas (1/1)
mot (36/36)
närarbetefinska (1/1)
sukupuolitautien (1/1)
orsakat (4/4)
bedömningsskalan (1/1)
stred (2/2)
värkjouren (1/1)
värnplikt (1/1)
könumret (1/1)
handpenning (1/1)
skapandet (1/1)
Mina (4/4)
köpingen (1/1)
preventivrådgivningen (1/1)
vård (57/57)
erityisammattitutkinto (1/1)
låter (1/1)
arbetarskyddet (2/2)
behörighet (4/4)
tulkki (1/1)
familjepension (5/5)
täydennyskoulutus (1/1)
flyktingorganisation (2/2)
fundera (8/8)
intressebevakningsorganisation (3/3)
följ (1/1)
förmånlig (2/2)
privatläkare (4/4)
måltidstjänst (1/1)
gjorts (1/1)
UNHCR:s (3/3)
pensionstagare (3/3)
sopsäck (1/1)
insikt (1/1)
bostadssökandet (1/1)
faktor (1/1)
skyddsåldersgränsen (1/1)
hormonella (2/2)
redskapet (1/1)
toalettstolen (1/1)
kunnig (1/1)
transportera (1/1)
IB (1/1)
middag (1/1)
rörelsenedsättning (2/2)
avbrott (9/9)
telefonservicefinska (1/1)
grenförbunden (1/1)
näyttötutkinto (4/4)
någonting (2/2)
påverkanfinska (1/1)
skolorna (5/5)
yrkeshögskolanfinska (2/2)
flyg (3/3)
barnlöshetsklinik (1/1)
lämningar (1/1)
orter (20/20)
II (1/1)
auttamisjärjestelmä (1/1)
sjukvård (8/8)
radhuslägenheter (1/1)
avlopp (2/2)
barnskyddslagenfinska (1/1)
R (1/1)
-flickor (1/1)
lämnar (12/12)
kuvataidekoulu (1/1)
pensionsskyddet (2/2)
arbetsuppgifter (8/8)
nätverk (9/9)
förbjuden (2/2)
lukio (4/4)
turvallisuusvirasto (1/1)
apoteken (1/1)
beredskap (1/1)
barnatillsyningsmannen (10/10)
arbete (78/82) Arbete (4)
Jesusbarnet (1/1)
hushållets (1/1)
bilagor (6/6)
bestyren (1/1)
flaggan (2/2)
jobbsökningscoachning (1/1)
nyheter (2/2)
dolda (1/1)
förvärvsarbeta (3/3)
barnskötare (3/3)
Erasmus (2/2)
social (12/12)
applikationsbutiken (1/1)
skuldrådgivarefinska (1/1)
dagvårdsstart (1/1)
sevärdheter (1/1)
Andelsbanken (1/1)
avgiftsbelagd (12/12)
avsedd (39/39)
hemmetfinska (1/1)
företagsverksamheten (9/9)
forskning (5/5)
tvärvetenskapliga (1/1)
saknar (6/6)
parten (3/3)
identifiera (2/2)
familjelivet (1/1)
flyttservice (1/1)
invånarnas (1/1)
tillsätter (1/1)
intill (3/3)
klubbarfinska (1/1)
hälft (1/1)
beskickningarna (1/1)
arbetsplatssajtfinska (1/1)
yrkeshögskoleexamenfinska (1/1)
kärnkraftverksprojekt (1/1)
Nuorten (3/3)
nioårig (1/1)
livshotande (2/2)
grundat (2/2)
medlemskommunernas (1/1)
rörande (3/3)
förmedlare (1/1)
säkerheter (1/1)
familjeåterföreningen (1/1)
undervisningsgrupper (1/1)
huvudsak (3/3)
trappuppgången (1/1)
linjekartor (1/1)
tillhörighet (3/3)
polisstation (1/1)
kapitalinkomsten (1/1)
stödåtgärder (1/1)
vuxengymnasier (2/2)
utmattade (1/1)
centralmuseetfinska (1/1)
intressebevakare (1/1)
emellertid (9/9)
tabletdator (1/1)
denne (3/3)
legaliserade (1/1)
uppdateringen (1/1)
personbeteckningar (1/1)
engelskspråkigt (1/1)
minderåriga (7/7)
el (3/3)
terveydenhoitaja (2/2)
tutkinta (1/1)
oroliga (1/1)
medborgarorganisation (1/1)
informera (1/1)
grundutbildning (2/2)
regiontrafiken (1/1)
vårens (1/1)
läkarhjälp (1/1)
stressyndrom (1/1)
vattentrafiken (1/1)
maistraatti (16/16)
informationfinska (1/1)
upptäckt (1/1)
handläggningen (2/2)
föreslog (1/1)
textinnehåll (1/1)
bildkonstskolor (1/1)
återflyttningfinska (1/1)
nödinkvartering (2/2)
av (1120/1120)
garantipension (2/2)
tis. (1/1)
statlig (1/1)
upptäcks (2/2)
bruttoinkomster (1/1)
hemskickad (1/1)
Flickornas (2/2)
döden (1/1)
Apostilleavtaletengelska (1/1)
pensionärer (4/4)
familjemedlemmarnas (2/2)
föreningens (3/3)
började (6/6)
r.f. (4/4)
förskolanfinska (1/1)
omedelbar (5/5)
öppenvården (1/1)
bostadens (9/9)
fart (1/1)
dygn (3/3)
samtalskostnad (1/1)
loven (1/1)
kortvarig (4/4)
jämnt (5/5)
anspråkslöshet (1/1)
kallt (3/3)
arbetsavtalfinska (1/1)
offentligt (7/7)
prövningsbaserat (1/1)
skryter (1/1)
omsorg (2/2)
bereda (1/1)
dags (1/1)
upphovsrätt (6/6)
eller (1301/1301)
konfidentiell (1/1)
TV:n (1/1)
täcka (5/5)
nöjd (1/1)
Oy (9/9)
Varias (1/1)
studiematerial (1/1)
Villa (1/1)
Medborgarrådgivning (1/1)
skolelevers (1/1)
vattenmätare (1/1)
högskolenivå (1/1)
gymnasieutbildningfinska (1/1)
turkiska (15/15)
utgående (8/8)
födelseattester (3/3)
FPAfinska (1/1)
Begravningsbyråers (1/1)
psykoterapeut (1/1)
korrigera (1/1)
grupp (9/9)
obligatoriskt (3/3)
utgifter (5/5)
håller (11/11)
levnadskostnaderna (1/1)
dagvårdenfinska (1/1)
upphävande (1/1)
parterna (7/7)
granska (1/1)
turvakoti (4/6) Turvakoti (2)
arbetslöshetsdagpenning (2/2)
slutet (14/14)
dem (64/64)
avslagits (1/1)
arbetstagarefinska (1/1)
riksdagen (2/2)
fysioterapeut (1/1)
tidsbokningen (5/5)
ryskaryska (1/1)
startade (1/1)
bidra (2/2)
tulkkikeskus (1/1)
reser (5/5)
företagshälsovårdenfinska (1/1)
Martinus (1/1)
hav (1/1)
idrottsgrenar (3/3)
karaoke (1/1)
upphävs (2/2)
förarexamen (1/1)
feber (1/1)
läkarintyget (1/1)
bekänner (2/2)
ritualer (1/1)
fastställer (2/2)
