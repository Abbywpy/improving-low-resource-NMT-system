då upphörde Saul att förfölja David och drog mot filistéerna . Därav fick det stället namnet Sela @-@ Hammalekot .
men själva kunna vi icke åt dem giva hustrur av våra döttrar , ty Israels barn hava svurit och sagt : Förbannad vare den som giver en hustru åt Benjamin &quot; .
då gingo de fem männen vidare och kommo till Lais ; och de sågo huru folket därinne bodde i trygghet , på sidoniernas sätt , stilla och trygga , och att ingen gjorde någon skada i landet genom att tillvälla sig makten ; och de bodde långt ifrån sidonierna och hade intet att skaffa med andra människor .
Filippus skyndade fram och hörde att han läste profeten Esaias . då frågade han : &quot; förstår du vad du läser ? &quot;
jag vill lyfta Mina händer upp till dina bud , ty de äro mig kära , och jag vill begrunda dina stadgar .
de omringa mig , ja , de omringa mig , men i HERRENS namn skall jag förgöra dem .
och var och en av dem förde med sig skänker : föremål av silver och av guld , kläder , vapen , välluktande kryddor , hästar och mulåsnor . så skedde år efter år .
då berövas de ogudaktiga sitt ljus , och den arm som lyftes för högt brytes sönder .
den rättfärdiges förvärv bliver honom till liv ; den ogudaktiges vinning bliver honom till synd .
men Jojada blev gammal och mätt på att leva och dog så ; ett hundra trettio år gammal var han vid sin död .
och de gjorde så och läto dem alla lägga sig ned .
och när de så , under sin flykt för Israel , hade kommit till den sluttning som går ned från Bet @-@ Horon , lät HERREN stora stenar falla över dem från himmelen , hela vägen ända till Aseka , så att de blevo dödade ; de som dödades genom hagelstenarna voro till och med flera än de som Israels barn dräpte med svärd .
och Jesus växte till i ålder och vishet och nåd inför Gud och människor .
och det fick en mun sig given , som talade stora ord och vad hädiskt var , och det fick makt att så göra under fyrtiotvå månader .
de skulle nämligen fråga prästerna i HERREN Sebaots hus och profeterna sålunda : &quot; skola vi framgent hålla gråtodag och späka oss i femte månaden , såsom vi hava gjort nu i så många år ? &quot;
den fostrar oss till att avsäga oss all ogudaktighet och alla världsliga begärelser , och till att leva tuktigt och rättfärdigt och gudfruktigt i den tidsålder som nu är ,
och konungen ropade med hög röst och befallde att man skulle hämta besvärjarna , kaldéerna ock stjärntydarna . och konungen lät säga så till de vise i Babel : &quot; Vemhelst som kan läsa denna skrift och meddela mig dess uttydning , han skall bliva klädd i purpur , och den gyllene kedjan skall hängas om hans hals , och han skall bliva den tredje herren i riket &quot; .
och när man hade offrat brännoffret , sade Jehu till drabanterna och kämparna : &quot; Gån in och slån ned dem ; låten ingen komma ut &quot; . och de slogo dem med svärdsegg , och drabanterna och kämparna kastade undan deras kroppar . därefter gingo de in i det Inre av Baals tempel
och det skall ske på den tiden att jag skall göra Jerusalem till en lyftesten för alla folk ; var och en som försöker lyfta den skall illa sarga sig därpå . och alla jordens folk skola församla sig mot det .
och prästen skall av offret taga en handfull , det som utgör själva altaroffret , och förbränna det på altaret ; därefter skall han giva kvinnan vattnet att dricka .
Hälsen alla bröderna med en helig kyss .
vidare Ajalon med dess utmarker och Gat @-@ Rimmon med dess utmarker ;
och ändå säga de av Israels hus : &quot; Herrens väg är icke alltid densamma &quot; ! skulle verkligen Mina vägar icke alltid vara desamma , I av Israels hus ? är det icke fastmer eder väg som icke alltid är densamma ?
men kommen ihåg , I Mina älskade , vad som har blivit förutsagt av vår Herres , Jesu Kristi , apostlar ,
till de andra åter säger jag själv , icke Herren : om någon som hör till bröderna har en hustru som icke är troende , och denna är villig att leva tillsammans med honom , så må han icke förskjuta henne .
vi vilja icke lämna eder , käre bröder , i okunnighet om huru det förhåller sig med dem som avsomna , för att I icke skolen sörja såsom de andra , de som icke hava något hopp .
och i första månaden , på fjortonde dagen i månaden , är HERRENS påsk .
är en man som bedrager sin nästa och sedan säger : &quot; jag gjorde det ju på skämt &quot; .
nej , hellre vill jag nu bliva kvävd , hellre dö än vara blott knotor !
han som icke har skonat sin egen Son , utan utgivit honom för oss alla , huru skulle han kunna annat än också skänka oss allt med honom ?
så skall det gå den glada staden , som satt så trygg , och som sade i sitt hjärta : &quot; jag och ingen annan ! &quot; Huru har den icke blivit en ödemark , en lägerstad för vilda djur ! alla som gå där fram skola vissla åt den och slå ihop händerna .
såsom HERREN hade bjudit Mose så hade Israels barn i alla stycken gjort allt arbete .
de hava öron och lyssna icke till , och ingen ande är i deras mun .
med honom är en arm av kött , men med oss är HERREN , vår Gud , och han skall hjälpa oss och föra våra krig . och folket tryggade sig vid Hiskias , Juda konungs , ord .
men det skall ske att var och en som åkallar HERRENS namn han skall varda frälst . Ty på Sions berg och i Jerusalem skall finnas en räddad skara , såsom HERREN har sagt ; och till de undsluppna skola höra de som HERREN kallar .
då räckte Aron ut sin hand över Egyptens vatten , och paddor stego upp och övertäckte Egyptens land .
så gick Åklagaren bort ifrån HERRENS ansikte och slog Job med svåra bulnader , ifrån fotbladet ända till hjässan .
och jag betraktade det och gav akt därpå ; då fick jag däri se fyrfota djur , sådana som leva på jorden , tama och vilda , så ock krälande djur och himmelens fåglar .
en annan sträcka sattes i stånd av Malkia , Harims son , och av Hassub , Pahat @-@ Moabs son , och därjämte Ugnstornet .
därefter sade han : &quot; tag pilarna &quot; . och när han hade tagit dem , sade han till Israels konung : &quot; slå på jorden &quot; . då slog han tre gånger och sedan höll han upp .
femton alnar högt steg vattnet över bergen , så att de övertäcktes .
i två hela år bodde han sedan kvar i en bostad som han själv hade hyrt . och alla som kommo till honom tog han emot ;
hos honom är väldighet och förskräckande makt , hos honom , som skapar frid i sina himlars höjd .
och därvid kommer det icke an på om någon är grek eller jude , omskuren eller oomskuren , barbar eller skyt , träl eller fri ; nej , Kristus är allt och i alla .
sedan gick allt folket hem , var och en till sitt ; men David vände om för att hälsa sitt husfolk .
sina gärningars kraft har han gjort kunnig för sitt folk , i det han gav dem hedningarnas arvedel .
och han skall döma mellan hednafolken och skipa rätt åt många folk . då skola de smida sina svärd till plogbillar och sina spjut till vingårdsknivar . Folken skola ej mer lyfta svärd mot varandra och icke mer lära sig att strida .
fursten Dison , fursten Eser , fursten Disan . dessa voro horéernas stamfurstar i Seirs land , var furste för sig .
när jag vill hela Israel , då uppenbarar sig Efraims missgärning och Samariens ondska . Ty de öva falskhet , tjuvar göra inbrott , rövarskaror plundra på vägarna .
och Israel kom till Egypten , Jakob blev en gäst i Hams land .
då alltså Edom icke tillstadde Israel att tåga genom sitt område , vek Israel av och gick undan för honom .
Onda andar blevo ock utdrivna ur många , och de ropade därvid och sade : &quot; du är Guds Son &quot; . men han tilltalade dem strängt och tillsade dem att icke säga något , eftersom de visste att han var Messias .
Ty jag är HERREN , som har fört eder upp ur Egyptens land , för att jag skall vara eder Gud . så skolen I nu vara heliga , ty jag är helig .
och jag skall sätta dem till att förrätta tjänsten i huset vid allt tjänararbete där , allt som där skall utföras .
av fäkreatur sjuttiotvå tusen ,
begär av mig , så skall jag giva dig hedningarna till arvedel och jordens ändar till egendom .
om någon icke förbliver i mig , så kastas han ut såsom en avbruten gren och förtorkas ; och man samlar tillhopa sådana grenar och kastar dem i elden , och de brännas upp .
och städerna Sodom och Gomorra lade han i aska och dömde dem till att omstörtas ; han gjorde dem så till ett varnande exempel för kommande tiders ogudaktiga människor .
då han nu vandrade utmed Galileiska sjön , fick han se två bröder , Simon , som kallas Petrus , och Andreas , hans broder , kasta ut nät i sjön , ty de voro fiskare .
Sannerligen säger jag eder : den stund kommer , jag , den är redan inne , så de döda skola höra Guds Sons röst , och de som höra den skola bliva levande .
var och en som hatar sin broder , han är en mandråpare ; och I veten att ingen mandråpare har evigt liv förblivande i sig .
men i stället hängåven I eder åt fröjd och glädje ; I dödaden oxar och slaktaden får , I åten kött och drucken vin , I saden : &quot; Låtom oss äta och dricka , ty i morgon måste vi dö &quot; .
och vilddjuret , som jag såg , liknade en panter , men det hade fötter såsom en björn och gap såsom ett lejon . och draken gav det sin makt och sin tron och gav det stor myndighet .
i andra raden en karbunkel , en safir och en kalcedon ;
om du stötte den oförnuftige mortel med en stöt , bland grynen , så skulle hans oförnuft ändå gå ur honom .
och det vart afton , och det vart morgon , den femte dagen .
och denna stadga skall du hålla på bestämd tid , år efter år .
sedan de hade ätit sig mätta , lättade de skeppet genom att kasta vetelasten i havet .
detta blev en orsak till synd ; folket gick ända till Dan för att träda fram inför den ena av dem .
HERREN är rättfärdig därinne , han gör intet orätt. var morgon låter han sin rätt gå fram i ljuset , den utebliver aldrig ; men de orättfärdiga veta icke av någon skam .
om du ser att den fattige förtryckes , och att rätt och rättfärdighet våldföres i landet , så förundra dig icke däröver ; ty på den höge vaktar en högre , och andra ännu högre vakta på dem båda .
Noa , Sem , Ham och Jafet .
se , detta står upptecknat inför Mina ögon ; jag skall icke tiga , förrän jag har givit vedergällning , ja , vedergällning i deras sköte ,
alltså , att han som förlänade eder Anden och utförde kraftgärningar bland eder gjorde detta , kom det sig av laggärningar eller därav att I lyssnaden i tro ,
men hennes handelsförvärv och vad hon får såsom skökolön skall vara helgat åt HERREN ; det skall icke läggas upp och icke gömmas , utan de som bo inför HERRENS ansikte skola av hennes handelsförvärv hava mat till fyllest och präktiga kläder .
i den församling som fanns i Antiokia verkade nu såsom profeter och lärare Barnabas och Simeon , som kallades Niger , och Lucius från Cyrene , så ock Manaen , landsfursten Herodes &apos; fosterbroder , och Saulus .
Ty HERREN Gud är sol och sköld ; HERREN giver nåd och ära ; han vägrar icke dem något gott , som vandra i ostrafflighet .
se , dagar skola komma , säger HERREN , då jag skall låta en rättfärdig telning uppstå åt David . han skall regera såsom konung och hava framgång , och han skall skaffa rätt och rättfärdighet på jorden .
då bugade sig Bat @-@ Seba , med ansiktet mot jorden , och föll ned för konungen och sade : &quot; må min herre , konung David , leva evinnerligen ! &quot;
och jag skall göra dem till ett enda folk i landet , på Israels berg ; en och samma konung skola de alla hava ; de skola icke mer vara två folk och icke mer vara delade i två riken .
för kehatiternas släkter föll lotten ut så , att bland dessa leviter prästen Arons söner genom lotten fingo ur Juda stam , ur simeoniternas stam och ur Benjamins stam tretton städer .
och alla flyktingar ur alla hans härskaror skola falla för svärd , och om några bliva räddade , så skola de varda förströdda åt alla väderstreck . och I skolen förnimma att jag , HERREN , har talat .
Ty konungen hade en egen Tarsisflotta på havet jämte Hirams flotta ; en gång vart tredje år kom Tarsisflottan hem och förde med sig guld och silver , elfenben , apor och påfåglar .
Låt min muns frivilliga offer behaga dig , HERRE , och lär mig dina rätter .
det ena som det andra har jag sett under Mina fåfängliga dagar : mången rättfärdig som har förgåtts i sin rättfärdighet , och mången orättfärdig som länge har fått leva i sin ondska .
dock , huru skulle det kunna få ro , då det är HERRENS bud det utför ? mot Askelon , mot Kustlandet vid havet , mot dem har han bestämt det .
då sade han till sina tjänare : &quot; i sen att Joab där har ett åkerstycke vid sidan av mitt , och på det har han korn ; gån nu dit och tänden eld därpå &quot; . så tände då Absaloms tjänare eld på åkerstycket .
och närmast Simeons område skall Isaskar hava en lott , från östra sidan till västra .
och Saul talade med sin son Jonatan och med alla sina tjänare om att döda David ; men Sauls son Jonatan var David mycket tillgiven .
den som tror och bliver döpt , han skall bliva frälst ; men den som icke tror , han skall bliva fördömd .
och min ande fröjdar sig i Gud , min Frälsare .
så äro vi då alltid vid gott mod . vi veta väl att vi äro borta ifrån Herren , så länge vi äro hemma i kroppen ;
då gick han åstad och begynte förkunna i Dekapolis huru stora ting Jesus hade gjort med honom ; och alla förundrade sig .
och hela Juda gladde sig över eden ; ty de hade svurit den av allt sitt hjärta , och de sökte HERREN med hela sin vilja , och han lät sig finnas av dem , och han lät dem få ro på alla sidor .
så må du veta : när profeten talar i HERRENS namn , och det som han har talat icke sker och icke inträffar , då är detta något som HERREN icke har talat ; i förmätenhet har då profeten talat det ; du skall icke frukta för honom &quot; .
sedan fick jag i min syn höra en örn , som flög fram uppe i himlarymden , ropa med hög röst : &quot; Ve , ve , ve över jordens inbyggare , när de tre övriga änglar , som skola stöta i basun , låta sina basuner ljuda ! &quot;
jag skyndar mig och dröjer icke att hålla dina bud .
hos dig må icke finnas någon som låter sin son eller dotter gå genom eld , eller som befattar sig med trolldom eller teckentydning eller svartkonst eller häxeri ,
och varen framför allt uthålliga i eder Kärlek till varandra , ty &quot; kärleken överskyler en myckenhet av synder &quot; .
och såsom han uttydde för oss , så gick det . jag blev åter insatt på min plats , och den andre blev upphängd &quot; .
såsom ditt namn , o Gud , så når ock ditt lov intill jordens ändar ; din högra hand är full av rättfärdighet .
och må nu icke mitt blod falla på jorden fjärran ifrån HERRENS ansikte , då Israels konung har dragit ut för att söka efter en enda liten loppa , såsom man jagar rapphöns på bergen &quot; .
av invånarna i Bet @-@ Semes blevo ock många slagna , därför att de hade sett på HERRENS ark ; han slog sjuttio man bland folket , femtio tusen man . och folket sörjde däröver att HERREN hade slagit så många bland folket .
han kan icke undslippa mörkret ; hans telningar skola förtorka av hetta , och själv skall han förgås genom Guds muns anda .
och detta är lagen om spisoffret : Arons söner skola bära fram det inför HERRENS ansikte , till altaret .
och sade : &quot; om jag har funnit nåd för dina ögon , Herre , så må Herren gå med oss . Ty väl är det ett hårdnackat folk , men du vill ju förlåta oss vår missgärning och synd och taga oss till din arvedel &quot; .
och så skall över eder komma allt rättfärdigt blod som är utgjutet på jorden , ända ifrån den rättfärdige Abels blod intill Sakarias &apos; , Barakias &apos; sons blod , hans som I dräpten mellan templet och altaret .
se , jag skall sända en ängel framför dig , som skall bevara dig på vägen och föra dig till den plats som jag har utsett .
och det skall ske i kommande dagar att det berg där HERRENS hus är skall stå där fast grundat och vara det yppersta ibland bergen och upphöjt över andra höjder ; och alla hednafolk skola strömma dit ,
då stampade hästarnas hovar , när deras tappra ryttare jagade framåt , framåt .
redan för länge sedan , redan då Saul ännu var konung , var det du som var ledare och anförare för Israel . och till dig har HERREN , din Gud , sagt : du skall vara en herde för mitt folk Israel , ja , du skall vara en furste över mitt folk Israel &quot; .
vi tacka dig , o Gud , vi tacka dig . ditt namn är oss nära ; man förtäljer dina under .
därefter begav han sig till en stad som hette Nain ; och med honom gingo hans lärjungar och mycket folk .
Mose svarade : &quot; du har talat rätt ; jag skall icke vidare komma inför ditt ansikte &quot; .
han som var till i Guds @-@ skepnad , men icke räknade jämlikheten med Gud såsom ett byte ,
men du , människobarn , hör nu vad jag talar till dig ; var icke gensträvig såsom detta gensträviga släkte . öppna din mun och ät vad jag giver dig &quot; .
och han gav tecken åt dem med handen att de skulle tiga , och förtäljde för dem huru Herren hade fört honom ut ur fängelset . och han tillade : &quot; Låten Jakob och de andra bröderna få veta detta &quot; . sedan gick han därifrån och begav sig till en annan ort .
Blevo vi icke av honom aktade såsom främlingar , när han sålde oss ? sedan har han ju ock förtärt vad han fick i betalning för oss .
sedan vände de båda männen tillbaka och kommo ned från bergsbygden och gingo över floden och kommo så till Josua , Nuns son ; och de förtäljde för honom allt vad som hade vederfarits dem .
och man förde fram sju tjurar , sju vädurar och sju lamm , så ock sju bockar till syndoffer för riket och för helgedomen och för Juda ; och han befallde Arons söner , prästerna , att offra detta på HERRENS altare .
Konung Salomo offrade såsom slaktoffer tjugutvå tusen tjurar och ett hundra tjugu tusen av småboskapen . så invigdes Guds hus av konungen och allt folket .
en uppfostrare för oförståndiga , en lärare för enfaldiga , eftersom du i lagen har uttrycket för kunskapen och sanningen .
här gäller det för de heliga att hava ståndaktighet , för dem som hålla Guds bud och bevara tron på Jesus &quot; .
jag skall låta strömmar rinna upp på höjderna och källor i dalarna ; jag skall göra öknen till en vattenrik sjö och torrt land till källsprång .
och i Manasses , Efraims och Simeons städer ända till Naftali genomsökte han överallt husen .
om han ville uppenbara dig sin visdoms lönnligheter , huru han äger förstånd , ja , i dubbelt mått , då insåge du att Gud , dig till förmån , har lämnat åt glömskan en del av din missgärning .
då sprutade ormen ur sitt gap vatten efter kvinnan såsom en ström , för att strömmen skulle bortföra henne .
så se nu till ; ty HERREN har utvalt dig att bygga ett hus till helgedomen . var frimodig och gå till verket &quot; .
och ljusstaken var gjord på följande sätt : den var av guld i drivet arbete ; också dess fotställning och blommorna därpå voro i drivet arbete . efter det mönster som HERREN hade visat Mose hade denne låtit göra ljusstaken .
men profeten Natan , Benaja , hjältarna och sin broder Salomo inbjöd han icke .
vidare berättade sekreteraren Safan för konungen och sade : &quot; Prästen Hilkia har givit mig en bok &quot; . och Safan föreläste den för konungen .
dessa skaffade sig moabitiska hustrur ; den ena hette Orpa och den andra Rut .
vilka hava vågat sina liv för vår Herres , Jesu Kristi , namns skull .
jag kallade på Mina vänner , men de bedrogo mig . Mina präster och Mina äldste förgingos i staden , medan de tiggde sig mat för att stilla sin hunger .
Kina , Dimona , Adada ,
och HERREN , din Gud , skall förjaga dessa hedningar för dig , men blott småningom . du skall icke med hast få förgöra dem , på det att vilddjuren icke må föröka sig till din skada .
gick vidare söder om Skorpionhöjden och fram till sin , drog sig så upp söder om Kades @-@ Barnea , gick därefter framom Hesron och drog sig upp till Addar samt böjde sig sedan mot Karka .
och Josef fann nåd för hans ögon och fick betjäna honom . och han satte honom över sitt hus , och allt vad han ägde lämnade han i hans vård .
och om han ser ett tåg , ryttare par efter par , ett tåg av åsnor , ett tåg av kameler , då må han giva akt , noga giva akt &quot; .
ty jag säger eder att jag icke mer skall fira denna högtid , förrän den kommer till fullbordan i Guds rike &quot; .
då svarade han honom : &quot; Välan , jag skall ock häri göra dig till viljes ; jag skall icke omstörta den stad som du talar om .
sådan var den dröm som jag , konung Nebukadnessar , hade . och du , Beltesassar , må nu säga uttydningen ; ty ingen av de vise i mitt rike kan säga mig uttydningen , men du kan det väl , ty heliga gudars ande är i dig &quot; .
kvinnor funnos som fingo igen sina döda genom deras uppståndelse . andra läto sig läggas på sträckbänk och ville icke taga emot någon befrielse , i hopp om en så mycket bättre uppståndelse .
men i konung Joas &apos; tjugutredje regeringsår hade prästerna ännu icke satt i stånd vad som var förfallet på huset .
och jag skall låta din säd bliva såsom stoftet på jorden ; kan någon räkna stoftet på jorden , så skall ock din säd kunna räknas .
då upptändes Balaks vrede mot Bileam , och han slog ihop händerna . och Balak sade till Bileam : &quot; till att förbanna Mina fiender kallade jag dig hit , och se , du har i stället nu tre gånger välsignat dem .
och han sover , och han vaknar , och nätter och dagar gå , och säden skjuter upp och växer i höjden , han vet själv icke huru .
om en man än finge hundra barn och finge leva i många år , ja , om hans livsdagar bleve än så många , men hans själ icke finge njuta sig mätt av hans goda , och om han så bleve utan begravning , då säger jag : lyckligare än han är ett ofullgånget foster .
en livets källa är förståndet för den som äger det , men oförnuftet är de oförnuftigas tuktan .
och färdades genom Syrien och Cilicien och styrkte församlingarna .
och var och en av eder må taga sitt fyrfat och lägga rökelse därpå , och sedan bära sitt fyrfat fram inför HERRENS ansikte , två hundra femtio fyrfat ; du själv och Aron mån ock taga var sitt fyrfat &quot; .
och David sade till honom : &quot; ditt blod komme över ditt huvud , ty din egen mun har vittnat mot dig , i det att du sade : &apos; jag har dödat HERRENS smorde . &apos; &quot;
och amoréerna förmådde hålla sig kvar i har @-@ Heres , Ajalon och Saalbim ; men Josefs barns hand blev tung över dem , så att de blevo arbetspliktiga under dessa .
sen icke därpå att jag är så svart , att solen har bränt mig så . min moders söner blevo vreda på mig och satte mig till vingårdsvakterska ; min egen vingård kunde jag icke vakta .
Böjen edra öron hit och kommen till mig ; hören , så får eder själ leva . jag vill sluta med eder ett evigt Förbund : att I skolen undfå all den trofasta nåd jag har lovat David .
dina präster vare klädda i rättfärdighet , och dina fromma juble .
och Mose och Aron gjorde alla dessa under inför Farao ; men HERREN förstockade Faraos hjärta , så att han icke släppte Israels barn ut ur sitt land .
och när I kommen in i någon stad där man tager emot eder , så äten vad som sättes fram åt eder ,
Förbannen Meros , säger HERRENS ängel , ja , förbannen dess inbyggare , därför att de ej kommo HERREN till hjälp , HERREN till hjälp bland hjältarna .
så sade nu Gud till Noa : &quot; detta skall vara tecknet till det Förbund som jag har upprättat mellan mig och allt kött på jorden &quot; .
men när Hiram från Tyrus begav sig ut för att bese de städer som Salomo hade givit honom , behagade de honom icke ,
så säger HERREN : se , jag skall uppväcka mot Babel och mot Leb @-@ Kamais inbyggare en fördärvares ande .
därför är jag villig att förkunna evangelium också för eder som bon i Rom .
och sedan Lemek hade fött Noa , levde han fem hundra nittiofem år och födde söner och döttrar .
Huru förvända ären I icke ! Skall då leret aktas lika med krukmakaren ? Skall verket säga om sin mästare : &quot; han har icke gjort mig &quot; ? eller skall bilden säga om honom som har format den : &quot; han förstår intet &quot; ?
jag skall låta min nitälskan gå över dig , så att de fara grymt fram mot dig ; de skola skära av dig näsa och öron , och de som bliva kvar av dig skola falla för svärd . man skall föra bort dina söner och döttrar , och vad som bliver kvar av dig skall förtäras av eld .
och somliga läto övertyga sig av det som han sade , men andra trodde icke .
Semaja , Jojarib , Jedaja ,
jag har ofta måst vara ute på resor ; jag har utstått faror på floder , faror bland rövare , faror genom landsmän , faror genom hedningar , faror i städer , faror i öknar , faror på havet , faror bland falska bröder --
när sabbaten hade gått till ända , i gryningen till första veckodagen , kommo Maria från Magdala och den andra Maria för att se graven .
vi hava funnit att denne är en fördärvlig man , som uppväcker strid bland alla judar i hela världen , och att han är en huvudman för nasaréernas parti .
varen såsom jag , som i alla stycken fogar mig efter alla och icke söker min egen nytta , utan de mångas , för att de skola bliva frälsta .
Amrams söner voro Aron och Mose . och Aron blev jämte sina söner för evärdlig tid avskild till att helgas såsom höghelig , till att för evärdlig tid antända rökelse inför HERREN och göra tjänst inför honom och välsigna i hans namn .
och framför vaktkamrarna var en avskrankning , som höll en aln ; en aln höll ock avskrankningen på motsatta sidan ; och var vaktkammare , på vardera sidan , höll sex alnar .
alltså , Mina älskade bröder , varen fasta , orubbliga , alltid överflödande i Herrens verk , eftersom I veten att edert arbete icke är fåfängt i Herren .
och när de nu förnummo vilken nåd som hade blivit mig given , räckte de mig och Barnabas handen till samarbete , både Jakob och Cefas och Johannes , de män som räknades för själva stödjepelarna ; vi skulle verka bland hedningarna , och de bland de omskurna .
och HERREN sade till honom : &quot; detta är det land som jag med ed har lovat åt Abraham . Isak och Jakob , i det jag sade : &apos; åt din säd skall jag giva det . &apos; jag har nu låtit dig se det med dina ögon , men ditin skall du icke komma &quot; .
när Baal @-@ Hanan , Akbors son , dog , blev Hadar konung efter honom ; och hans stad hette Pagu , och hans hustru hette Mehetabel , dotter till Matred , som var dotter till Me @-@ Sahab .
man bedriver styggelse , var och en med sin nästas hustru ; ja , man orenar i skändlighet sin sons hustru ; man kränker hos dig sin syster , sin faders dotter .
och HERRENS ord kom till mig ; han sade : du människobarn , säg till dem :
Strömportarna måste öppna sig , och palatset försmälter av ångest .
utan den plats som HERREN , eder Gud , utväljer inom någon av edra stammar till att där fästa sitt namn , denna boning skolen I söka och dit skall du gå .
ja , är det icke så med mitt hus inför Gud ? han har ju upprättat med mig ett evigt Förbund , i allo stadgat och betryggat . ja , visst skall han låta all frälsning och glädje växa upp åt mig .
Veten I då icke att de orättfärdiga icke skola få Guds rike till arvedel ? Faren icke vilse . varken otuktiga människor eller avgudadyrkare eller äktenskapsbrytare , varken de som låta bruka sig till synd mot naturen eller de som själva öva sådan synd ,
och han lät leviterna ställa upp sig till tjänstgöring i HERRENS hus med cymbaler , psaltare och harpor , såsom David och Gad , konungens siare , och profeten Natan hade bjudit ; ty budet härom var givet av HERREN genom hans profeter .
i de synderna vandraden också I förut , då I ännu haden edert liv i dem .
Konungen frågade honom &quot; Var är han ? &quot; Siba svarade konungen : &quot; han är nu i Makirs , Ammiels sons , hus i Lo @-@ Debar &quot; .
och härar , utsända av honom , skola komma och oskära helgedomens fäste och avskaffa det dagliga offret och ställa upp förödelsens styggelse .
här är icke jude eller grek , här är icke träl eller fri , här är icke man och kvinna : alla ären I ett i Kristus Jesus .
Kraftverkningarna äro mångahanda , men Gud är en och densamme , han som verkar allt i alla .
Lyft det sedan i deras åsyn upp på axeln och för bort det , när det har blivit alldeles mörkt ; och betäck ditt ansikte , så att du icke ser landet . Ty jag gör dig till ett tecken för Israels hus &quot; .
då sade jag till min herre : &apos; men om nu kvinnan icke vill följa med mig ? &apos;
allt såsom HERREN hade bjudit Mose ; och han mönstrade dem i Sinais öken .
hans huvud och hår var vitt såsom vit ull , såsom snö , och hans ögon voro såsom eldslågor .
men männen ville icke höra på honom ; då tog mannen sin bihustru och förde henne ut till dem . och de kände henne och hanterade henne skändligt hela natten ända till morgonen ; först när morgonrodnaden gick upp , läto de henne gå .
&quot; dessa voro de män från hövdingdömet , som drogo upp ur den landsflykt och fångenskap till vilken de hade blivit bortförda av Nebukadnessar , konungen i Babel , och som vände tillbaka till Jerusalem och till Juda , var och en till sin stad ,
Huru skall en yngling bevara sin väg obesmittad ? när han håller sig efter ditt ord .
den som har öra , han höre vad Anden säger till församlingarna &quot; .
och Faraos dotter kom ned till floden för att bada , och hennes tärnor gingo utmed floden . när hon nu fick se kistan i vassen , sände hon sin tjänarinna dit och lät hämta den till sig .
alla dessa höllo endräktigt ut i bön tillika med Maria , Jesu moder , och några andra kvinnor samt Jesu bröder .
och Saul och allt det folk som han hade hos sig församlade sig och drogo till stridsplatsen ; där fingo de se att den ene hade lyft sitt svärd mot den andre , så att en mycket stor förvirring hade uppstått .
Ty jag är viss om att varken död eller liv , varken änglar eller andefurstar , varken något som nu är eller något som skall komma ,
det må vara lärjungen nog , om det går honom såsom hans mästare , och tjänaren , om det går honom såsom hans herre . om de hava kallat husbonden för Beelsebul , huru mycket mer skola de icke så kalla hans husfolk !
därför säger HERREN så om Anatots män , dem som stå efter ditt liv och säga : &quot; Profetera icke i HERRENS namn , om du icke vill dö för vår hand &quot;
sedan trädde de fram till honom och sade : &quot; Hell dig , du judarnas konung ! &quot; och slogo honom på kinden .
åt denne inrett en stor kammare , där man förut plägade lägga in spisoffret , rökelsen och kärlen och den tionde av säd , vin och olja , som var bestämd åt leviterna , sångarna och dörrvaktarna , så ock offergärden åt prästerna .
ja , alla andra folk vandra vart och ett i sin guds namn , men vi vilja vandra i HERRENS , vår Guds , namn , alltid och evinnerligen .
när lärjungarna sågo detta , förundrade de sig och sade : &quot; Huru kunde fikonträdet så i hast förtorkas ? &quot;
och prästerna , Levi söner , skola träda fram , ty dem har HERREN , din Gud , utvalt till att göra tjänst inför honom och till att välsigna i HERRENS namn , och såsom de bestämma skola alla tvister och alla misshandlingsmål behandlas .
så ofta israeliterna hade sått , drogo midjaniterna , amalekiterna och österlänningarna upp emot dem
vid deras åsyn gripas folken av ångest , alla ansikten skifta färg .
och Aron var ett hundra tjugutre år gammal , när han dog på berget Hor .
i samma stund kommo några fariséer fram och sade till honom : &quot; Begiv dig åstad bort härifrån ; ty Herodes vill dräpa dig &quot; .
och han förde fram brännoffersväduren , och Aron och hans söner lade sina händer på vädurens huvud .
då trädde en av de skriftlärde fram , en som hade hört deras ordskifte och förstått att han hade svarat dem väl . denne frågade honom : &quot; vilket är det förnämsta av alla buden ? &quot;
eftersom I genom lögnaktigt tal haven gjort den rättfärdige försagd i hjärtat , honom som jag ingalunda ville plåga , men däremot haven styrkt den ogudaktiges mod , så att han icke vänder om från sin onda väg och räddar sitt liv ,
men alltsammans kommer från Gud , som har försonat oss med sig själv genom Kristus och givit åt oss försoningens ämbete .
men jag hämtade eder fader Abraham från andra sidan floden och lät honom vandra omkring i hela Kanaans land . och jag gjorde hans säd talrik ; jag gav honom Isak ,
och Farao blev förtörnad på sina två hovmän , överste munskänken och överste bagaren ,
då nu Jesus märkte att han hade svarat förståndigt , sade han till honom : &quot; du är icke långt ifrån Guds rike &quot; . sedan dristade sig ingen att vidare ställa någon fråga på honom .
och sade : &quot; Herre , min tjänare ligger därhemma lam och lider svårt &quot; .
då svarade allt folket med en mun och sade : &quot; allt vad HERREN har talat vilja vi göra &quot; . och Mose gick tillbaka till HERREN med folkets svar .
och om ditt offer är ett spisoffer som tillredes på plåt , så skall det vara av fint mjöl , begjutet med olja , osyrat .
och de talade inställsamt för honom med sin mun och skrymtade för honom med sin tunga .
om han vill bära fram ett brännoffer av fäkreaturen , så skall han därtill taga ett felfritt djur av hankön och föra det fram till uppenbarelsetältets ingång , för att han må bliva välbehaglig inför HERRENS ansikte .
på samma sätt hade han gjort för Esaus barn , som bo i Seir , i det han för dem förgjorde horéerna ; de fördrevo dem och bosatte sig i deras land , där de bo ännu i dag .
det bud som Jonadab , Rekabs son , gav sina barn , att de icke skulle dricka vin , det har blivit iakttaget , och ännu i dag dricka de icke vin , av hörsamhet mot sin faders bud . men själv har jag titt och ofta talat till eder , och I haven dock icke hörsammat mig .
och däri består kärleken , att vi vandra efter de bud han har givit . ja , detta är budet , att I skolen vandra i kärleken , enligt vad I haven hört från begynnelsen .
hon bliver ock agad genom plågor på sitt läger och genom ständig oro , allt intill benen .
Gören därför bättring och omvänden eder , så att edra synder bliva utplånade ,
men där var ock en annan stor örn med stora vingar och fjädrar i mängd ; och se , till denne böjde nu vinträdet längtansfullt sina grenar , och från platsen där det var planterat sträckte det sina rankor mot honom , för att han skulle vattna det .
jag vill höra vad Gud , HERREN , talar : se , han talar frid till sitt folk och till sina fromma ; må de blott icke vända åter till dårskap .
och hövding för gersoniternas stamfamilj var Eljasaf , Laels son .
Ty då hedningarna , som icke hava lag , av naturen göra vad lagen innehåller , så äro dessa , utan att hava lag , sig själv en lag ,
och konung David sade till hela församlingen : &quot; min son Salomo den ende som Gud har utvalt , är ung och späd , och arbetet är stort , ty denna borg är icke avsedd för en människa , utan för HERREN Gud .
då nu Jesus märkte att han hade svarat förståndigt , sade han till honom : &quot; du är icke långt ifrån Guds rike &quot; . sedan dristade sig ingen att vidare ställa någon fråga på honom .
och Mose och Aron och hans söner tvådde sedermera sina händer och fötter med vatten därur ;
&quot; Sannerligen , sannerligen säger jag eder : den som icke går in i fårahuset genom dörren , utan stiger in någon annan väg , han är en tjuv och en rövare .
den som ävlas att få vänner , han kommer i olycka ; men vänner finnas , mer trogna än en broder .
hans offergåva var ett silverfat , ett hundra trettio siklar i vikt , och en silverskål om sjuttio siklar , efter helgedomssikelns vikt , båda fulla med fint mjöl , begjutet med olja , till spisoffer ,
genom att höra på dem förökar den vise sin lärdom och förvärvar den förståndige rådklokhet .
och du , människobarn , profetera och såg : så säger Herren , HERREN om Ammons barn och om deras smädelser : Säg : ett svärd , ja , ett svärd är draget , det är fejat för att slakta för att varda mättat och för att blixtra ,
därför skall deras väg bliva för dem såsom en slipprig stig i mörkret , de skola på den stöta emot och falla . Ty jag vill låta olycka drabba dem , när deras hemsökelses är kommer , säger HERREN .
Låten båda slagen växa tillsammans intill skördetiden ; och när skördetiden är inne , vill jag säga till skördemännen : &apos; Samlen först tillhopa ogräset , och binden det i knippor till att brännas upp , och samlen sedan in vetet i min lada . &apos; &quot;
men de ropade till HERREN i sin nöd , och han frälste dem ur deras trångmål ;
det lilla som en rättfärdig har är bättre än många ogudaktigas stora håvor .
det är icke I som skolen tala , utan det är eder Faders Ande som skall tala i eder .
och HERREN bjöd oss att göra efter all dessa stadgar och att frukta HERREN , vår Gud , för att det alltid skulle gå oss väl , i det att han behölle oss vid liv , såsom ock hittills har skett .
och Gud välsignade dem ; Gud sade till dem : &quot; Varen fruktsamma och föröken eder , och uppfyllen jorden och läggen den under eder ; och råden över fiskarna i havet och över fåglarna under himmelen och över alla djur som röra sig på jorden &quot; .
dina heliga städer hava blivit en öken , Sion har blivit en öken , Jerusalem en ödemark .
och han lät oss komma hit och gav oss detta land , ett land som flyter av mjölk och honung .
om nu Satan driver ut Satan , så har han kommit i strid med sig själv . Huru kan då hans rike hava bestånd ?
så föllo av Benjamin aderton tusen man , allasammans tappert folk .
och vad du måste utbetala för det som härutöver behöves till din Guds hus , det må du låta utbetala ur konungens skattkammare .
Tjänen HERREN med glädje , kommen inför hans ansikte med fröjderop .
och ur korgen med de osyrade bröden , som stod inför HERRENS ansikte , tog han en osyrad kaka , en oljebrödskaka och en tunnkaka och lade detta på fettstyckena och det högra lårstycket .
och fönster funnos på den och på dess förhus runt omkring , likadana som de andra fönstren . den var femtio alnar lång och tjugufem alnar bred .
ja , klagoropen ljuda runtom i Moabs land ; till Eglaim når dess jämmer och till Beer @-@ Elim dess jämmer .
utan du skall gå till den plats som Herren , din Gud , utväljer till boning åt sitt namn , och där skall du slakta påskoffret om aftonen , när solen går ned den tid på dagen , då den drog ut ur Egypten .
Ty en annan grund kan ingen lägga , än den som är lagd , nämligen Jesus Kristus ;
och ingen annan rökelse mån I göra åt eder så sammansatt som denna skall vara . Helig skall den vara dig för HERREN .
och striden blev på den dagen allt häftigare , och Israels konung höll sig ända till aftonen upprätt i sin vagn , vänd mot araméerna ; men vid den tid då solen gick ned gav han upp andan .
Vaken , och bedjen att I icke mån komma i frestelse . Anden är villig , men köttet är svagt &quot; .
då svarade Jesus honom : &quot; Rävarna hava kulor , och himmelens fåglar hava nästen ; men Människosonen har ingen plats där han kan vila sitt huvud &quot; .
ett falskt vittne bliver icke ostraffat , och den som främjar lögn , han kommer icke undan .
Likväl sänder jag nu åstad dessa bröder , för att det som jag har sagt till eder berömmelse icke skall i denna del befinnas hava varit tomt tal . Ty , såsom jag förut har sagt , jag vill att I skolen vara redo .
Kallar jag på min tjänare , så svarar han icke ; ödmjukt måste jag bönfalla hos honom .
och över judarnas äldste vakade deras Guds öga , så att man lovade att icke lägga något hinder i vägen för dem , till dess saken hade kommit inför Darejaves ; sedan skulle man sända dem en skrivelse härom .
Konungen frågade : &quot; Finnes ingen kvar av Sauls hus , mot vilken jag kan bevisa barmhärtighet , såsom Gud är barmhärtig ? &quot; Siba svarade konungen : &quot; ännu finnes kvar en son till Jonatan , en som är ofärdig i fötterna &quot; .
han höll nämligen Kristi smälek för en större rikedom än Egyptens skatter , ty han hade sin blick riktad på lönen .
ty du vet att en sådan är förvänd och begår synd , ja , han har själv fällt domen över sig .
den som fruktar HERREN , han vandrar i redlighet , men den som föraktar honom , han går krokiga vägar .
Väduren som du såg , han med de två hornen , betyder Mediens och Persiens konungar .
där uppehöll han sig i tre månader . när han sedan tänkte avsegla därifrån till Syrien , beslöt han , eftersom judarna förehade något anslag mot honom , att göra återfärden genom Macedonien .
och överhovmästaren Eljakim och sekreteraren Sebna och de äldste bland prästerna sände han , höljda i sorgdräkt , till profeten Jesaja , Amos &apos; son .
och du skall göra femtio häktor av guld och foga tillhopa våderna med varandra medelst häktorna , så att tabernaklet utgör ett helt .
och sade : &quot; så skolen I säga : &apos; hans lärjungar kommo om natten och stulo bort honom , medan vi sovo . &apos;
av den minste skola komma tusen , och av den ringaste skall bliva ett talrikt folk . jag är HERREN ; när tiden är inne , skall jag med hast fullborda detta .
och de bådo och sade : &quot; Herre , du som känner allas hjärtan , visa oss vilken av dessa två du har utvalt
bjöd han leviterna som buro HERRENS förbundsark och sade :
Gören därför bättring och omvänden eder , så att edra synder bliva utplånade ,
Ty väl är det fåfängt , då man vill fånga fåglar , att breda ut nätet i hela flockens åsyn .
och var och en som icke gör efter din Guds lag och konungens lag , över honom skall dom fällas med rättvisa , vare sig till död eller till landsförvisning eller till penningböter eller till fängelse &quot; .
ja , förstår du himmelens lagar , och ordnar du dess välde över jorden ?
men de stodo stilla , var och en på sin plats , runt omkring lägret . då begynte alla i lägret att löpa hit och dit och skria och fly .
må deras bord framför dem bliva till en snara och till ett giller , bäst de gå där säkra ;
det har blivit ditt fördärv , o Israel , att du satte dig upp mot mig som var din hjälp .
men Jonatan , Davids farbroder , var rådgivare ; han var en förståndig och skriftlärd man . Jehiel , Hakmonis son , var anställd hos konungens söner .
av Josefs barn : av Efraim : Elisama , Ammihuds son ; av Manasse : Gamliel , Pedasurs son ;
fick han fatt på en ung man , en av invånarna i Suckot , och utfrågade denne , och han måste skriva upp åt honom de överste i Suckot och de äldste där , sjuttiosju män .
och Hosea , Elas son , anstiftade en sammansvärjning mot Peka , Remaljas son , och slog honom till döds och blev så konung i hans ställe , i Jotams , Ussias sons , tjugonde regeringsår .
men kaldéernas här förföljde konungen , och de hunno upp honom på Jerikos hedmarker , sedan hela hans här hade övergivit honom och skingrat sig .
Ty var och en som beder , han får ; och den som söker , han finner ; och för den som klappar skall varda upplåtet .
du skall trolova dig med en kvinna , men en annan man skall sova hos henne ; du skall bygga ett hus , men icke få bo däri ; du skall plantera en vingård , men icke få skörda dess frukt .
om jag nu har anbefallt Titus , så mån I besinna att han är min medbroder och min medarbetare till edert bästa ; och om jag har skrivit om andra våra bröder , så mån I besinna att de äro församlingssändebud och Kristi ära .
eftersom du är så dyrbar i Mina ögon , så högt aktad och så älskad av mig , därför giver jag människor till lösen för dig och folk till lösen för ditt liv .
Mina sabbater skolen I hålla , och för min helgedom skolen I hava fruktan . jag är HERREN .
hedningarna åter hava fått prisa Gud för hans barmhärtighets skull . så är ock skrivet : &quot; Fördenskull vill jag prisa dig bland hedningarna och lovsjunga ditt namn &quot; .
ditt majestäts härlighet och ära vill jag begrunda och dina underfulla verk .
men somt föll i god jord , och det sköt upp och växte och gav frukt och bar trettiofalt och sextiofalt och hundrafalt &quot; .
men när han hörde detta , blev han djupt bedrövad , ty han var mycket rik .
vad orsak haven I till att bruka detta ordspråk i Israels land : &quot; Fäderna äta sura druvor , och barnens tänder bliva ömma därav &quot; ?
och Jakob flydde till Arams mark Israel tjänade för en kvinna , för en kvinnas skull vaktade han hjorden .
och han kom tillbaka till Juda och sade : &quot; jag har icke funnit henne ; därtill säger folket på orten att ingen tempeltärna har varit där &quot; .
det har varit för mig en stor glädje i Herren att I nu omsider haven kommit i en så god ställning , att I haven kunnat tänka på mitt bästa . dock , I tänkten nog också förut därpå , men I haden icke tillfälle att göra något .
Kus &apos; söner voro Seba , Havila , Sabta , Raema och Sabteka . Raemas söner voro Saba och Dedan .
Uppe på höjderna står hon , vid vägen , där stigarna mötas .
om någon icke vill omvända sig , så vässer han sitt svärd , sin båge spänner han och gör den redo ;
Esau sade till sin fader : &quot; har du då allenast den enda välsignelsen , min fader ? Välsigna också mig , min fader &quot; . och Esau brast ut i gråt .
HERREN är sitt folks starkhet , och ett frälsningens värn är han för sin smorde .
då han emellertid ville få säkert besked om varför Paulus anklagades av judarna , låt han dagen därefter taga av honom bojorna och bjöd översteprästerna och hela Stora rådet att komma tillsammans . sedan lät han föra Paulus ditned och ställde honom inför dem .
om en prästs dotter ohelgar sig genom skökolevnad , så ohelgar hon sin fader ; hon skall brännas upp i eld .
fattade hon honom i manteln och sade : &quot; Ligg hos mig &quot; . men han lämnade manteln i hennes hand och flydde och kom ut .
då sade han till honom : &quot; eftersom du icke har lyssnat till HERRENS röst , därför skall ett lejon slå ned dig , när du går ifrån mig &quot; . och när han gick sin väg ifrån honom , kom ett lejon emot honom och slog ned honom .
ej heller skall du i ditt hus hava två slags efa @-@ mått , ett större och ett mindre .
Folket , som stod där och hörde detta , sade då : &quot; det var ett tordön &quot; . andra sade : &quot; det var en ängel som talade med honom &quot; .
Sion hör det och gläder sig , och Juda döttrar fröjda sig för dina domars skull , HERRE .
här visade sig för Paulus i en syn om natten en macedonisk man , som stod där och bad honom och sade : &quot; far över till Macedonien och hjälp oss &quot; .
upp , alla I som ären törstiga , kommen hit och fån vatten ; och I som inga penningar haven , kommen hit och hämten säd och äten . ja , kommen hit och hämten säd utan penningar och för intet både vin och mjölk .
Tänk , min Gud på Tobia , ävensom Sanballat , efter dessa hans gärningar , så ock på profetissan Noadja och de andra profeterna som ville skrämma mig !
men jag har något litet emot dig : du har hos dig några som hålla fast vid Balaams lära , hans som lärde Balak huru han skulle lägga en stötesten för Israels barn , så att de skulle äta kött från avgudaoffer och bedriva otukt .
då nu Moses svärfader såg allt vad han hade att beställa med folket , sade han : &quot; vad är det allt du har att bestyra med folket ? varför sitter du här till doms ensam under det att allt folket måste stå omkring dig från morgonen ända till aftonen ? &quot;
för sångmästaren ; av Koras söner ; en psalm .
Ty deras vredes stora dag är kommen , och vem kan bestå ? &quot;
och Hiskia gick till vila hos sina fäder . och hans son Manasse blev konung efter honom .
och till Amasa skolen I säga : &apos; är du icke mitt kött och ben ? Gud straffe mig nu och framgent , om du icke för all din tid skall bliva härhövitsman hos mig i Joabs ställe . &apos; &quot;
så skall då Herren , HERREN Sebaot sända tärande sjukdom i hans feta kropp , och under hans härlighet skall brinna en brand likasom en brinnande eld .
Ty dessa lade alla dit av sitt överflöd , men hon lade dit av sitt armod allt vad hon hade , så mycket som fanns i hennes ägo &quot; .
och de fem män som hade varit åstad för att bespeja landet gingo upp och kommo ditin och togo den skurna gudabilden och efoden , så ock husgudarna och den gjutna gudabilden , under det att prästen stod vid ingången till porten jämte de sex hundra vapenomgjordade männen .
jag levde en gång utan lag ; men när budordet kom , fick synden liv ,
vi älska dem för sanningens skull , som förbliver i oss , och som skall vara med oss till evig tid .
detta är vad som stod i det brev som profeten Jeremia sände från Jerusalem till de äldste som ännu levde kvar i fångenskapen , och till prästerna och profeterna och allt folket , dem som Nebukadnessar hade fört bort ifrån Jerusalem till Babel ,
Förhuset var tjugu alnar lång och elva alnar brett , nämligen vid trappstegen på vilka man steg ditupp . och vid murpelarna stodo pelare , en på var sida .
när Hirams flotta hämtade guld från Ofir , hemförde också den från Ofir almugträ i stor myckenhet , ävensom ädla stenar .
Skära mig med isop , så att jag varder ren ; två mig , så att jag bliver vitare än snö .
Ty det ordet skulle fullbordas , som han hade sagt : &quot; av dem som du har givit mig har jag icke förlorat någon &quot; .
239400
en bihustru som han hade i Sikem födde honom ock en son ; denne gav han namnet Abimelek .
icke är jag väl ett hav eller ett havsvidunder , så att du måste sätta ut vakt mot mig ?
Låt varna dig , Jerusalem , så att min själ ej vänder sig ifrån dig , så att jag icke gör dig till en ödemark , till ett obebott land .
och Jesus talade till honom och sade : &quot; vad vill du att jag skall göra dig ? &quot; den blinde svarade honom : &quot; Rabbuni , låt mig få min syn &quot; .
Ben @-@ Geber i Ramot i Gilead ; han hade Manasses son Jairs byar , som ligga i Gilead ; han hade ock landsträckan Argob , som ligger i Basan , sextio stora städer med murar och kopparbommar ;
och du skall älska HERREN , din Gud , av allt ditt hjärta och av all din själ och av all din kraft .
och Jakob sade till sina fränder : &quot; Samlen tillhopa stenar &quot; . och de togo stenar och gjorde ett röse och höllo måltid där på röset .
om däremot någon är fast i sitt sinne och icke bindes av något nödtvång , utan kan följa sin egen vilja , och så i sitt sinne är besluten att låta sin ogifta dotter förbliva såsom hon är , då gör denne väl .
och den som skall renas skall två sina kläder och raka av allt sitt hår och bada sig i vatten , så bliver han ren och får sedan gå in i lägret . dock skall han stanna utanför sitt tält i sju dagar .
de svulster av guld som filistéerna gåvo såsom skuldoffer åt HERREN utgjorde : för Asdod en , för Gasa en , för Askelon en , för Gat en , för Ekron en .
och Johannes hade kläder av kamelhår och bar en lädergördel om sina länder och levde av gräshoppor och vildhonung .
Ställ dig i porten till HERRENS hus , och predika där detta ord och säg : Hören HERRENS ord , I alla av Juda , som gån in genom dessa portar för att tillbedja HERREN .
när Saul nu hade tagit konungadömet över Israel i besittning , förde han krig mot alla sina fiender runt omkring : mot Moab , mot Ammons barn , mot Edom , mot konungarna i Soba och mot filistéerna ; och vart han vände sig tuktade han dem .
och Josef dog , när han var ett hundra tio år gammal . och man balsamerade honom , och han lades i en kista , i Egypten .
aviterna gjorde sig en Nibhas och en Tartak , och sefarviterna brände upp sina barn i eld åt Adrammelek och Anammelek , Sefarvaims gudar .
de befästa sig i sitt onda uppsåt , de orda om huru de skola lägga ut snaror ; de säga : &quot; vem skulle se oss ? &quot;
varhelst någon oförvitlig man funnes , en enda kvinnas man , en som hade troende barn , vilka icke vore i vanrykte för oskickligt leverne eller vore uppstudsiga .
och den omfattade Kattat , Nahalal , Simron , Jidala och Bet @-@ Lehem -- tolv städer med deras byar .
Mjölk gav jag eder att dricka ; fast föda gav jag eder icke , ty det fördrogen I då ännu icke . ja , icke ens nu fördragen I det ,
därför säger Herren , HERREN så : eftersom edert tal är falskhet och edra syner äro lögn , se , därför skall jag komma över eder , säger Herren , HERREN .
och HERRENS tjänare Mose dog där i Moabs land , såsom HERREN hade sagt .
Ty ljusets frukt består i allt vad godhet och rättfärdighet och sanning är .
och när folket såg honom , lovade de likaledes sin gud och sade : &quot; Vår gud har givit vår fiende i vår hand honom som förödde vårt land och slog så många av oss ihjäl &quot; .
när de hörde detta , prisade de Gud . och de sade till honom : &quot; du ser , käre broder , huru många tusen judar det är som hava kommit till tro , och alla nitälska de för lagen .
Lottkastning gör en ände på trätor , den skiljer mellan mäktiga män .
Visserligen har allt detta fått namn om sig att vara &quot; vishet &quot; , eftersom däri ligger ett självvalt gudstjänstväsende och ett slags &quot; ödmjukhet &quot; och en kroppens späkning ; men ingalunda ligger däri &quot; en viss heder &quot; , det tjänar allenast till att nära det köttsliga sinnet .
då svarade Jakob och sade till Laban : &quot; jag fruktade för dig , ty jag tänkte att du skulle med våld taga dina döttrar ifrån mig .
då drog konung Joram ut från Samaria och mönstrade hela Israel .
HERREN är konung evinnerligen , din Gud , Sion , från släkte till släkte . Halleluja !
men staden med allt vad däri är skall givas till spillo åt HERREN ; allenast skökan Rahab skall få leva , jämte alla som äro inne i hennes hus , därför att hon gömde de utskickade som vi hade sänt åstad .
så många av Efraims stam som inmönstrades ; utgjorde fyrtio tusen fem hundra .
men över Davids hus och över Jerusalems invånare skall jag utgjuta en nådens och bönens ande , så att de se upp till mig , och se vem de hava stungit . och de skola hålla dödsklagan efter honom , såsom man håller dödsklagan efter ende sonen , och skola bittert sörja honom , såsom man sörjer sin förstfödde .
Åter talade Jesus till dem och sade : &quot; jag är världens ljus ; den som följer mig , han skall förvisso icke vandra i mörkret , utan skall hava livets ljus &quot; .
Tagen därför ifrån honom hans pund , och given det åt den som har de tio punden .
eller är Gud allenast judarnas Gud ? är han icke ock hedningarnas ? Jo , förvisso också hedningarnas ,
i världen var han , och genom honom hade världen blivit till , men världen ville icke veta av honom .
så låtom oss lära känna HERREN , ja , låtom oss fara efter att lära känna honom . hans uppgång är så viss som morgonrodnadens , och han skall komma över oss lik ett regn , lik ett vårregn , som vattnar jorden &quot; .
åt denne gav då Simon Petrus ett tecken och sade till honom : &quot; Säg vilken det är som han talar om &quot; .
så många av Naftali stam som inmönstrades , utgjorde femtiotre tusen fyra hundra .
Rök steg upp från hans näsa och förtärande eld från hans mun ; eldsglöd ljungade från honom .
inom sina förtryckares murar måste de bereda olja , de få trampa vinpressar och därvid lida törst .
och Abram blev av honom väl behandlad för hennes skull , så att han fick får , fäkreatur och åsnor , tjänare och tjänarinnor , åsninnor och kameler .
gåvor öppna väg för en människa och föra henne fram inför de store .
nej , I gören eder faders gärningar &quot; . de sade till honom : &quot; vi äro icke födda i äktenskapsbrott . vi hava Gud till fader och ingen annan &quot; .
och jag skall sätta dem till att förrätta tjänsten i huset vid allt tjänararbete där , allt som där skall utföras .
därför , om nu en profet profeterar om lycka , så kan man först då när den profetens ord går i fullbordan veta att han är en profet som HERREN i sanning har sänt &quot; .
och edra altaren skola varda förödda och edra solstoder sönderkrossade , och dem av eder , som bliva slagna , skall jag låta bliva kastade inför edra eländiga avgudar .
Mosa födde Binea . hans son var Rafa ; hans son var Eleasa ; hans son var Asel .
om någon ligger hos sin svärdotter , så skola de båda straffas med döden ; de hava bedrivit en vederstygglighet , blodskuld låder vid dem .
jag sade i mitt hjärta : &quot; se , jag har förvärvat mig stor vishet , och jag har förökat den , så att den övergår allas som före mig hava regerat över Jerusalem ; ja , vishet och insikt har mitt hjärta inhämtat i rikt mått &quot; .
men när Cefas kom till Antiokia , trädde jag öppet upp mot honom , ty han hade befunnits skyldig till en försyndelse .
då skall du överlämna åt HERREN allt det som öppnar moderlivet . allt som öppnar moderlivet av det som födes bland din boskap skall , om det är hankön , höra HERREN till .
så att markens djur skola ära mig , schakaler och strutsar , därför att jag låter vatten flyta i öknen , strömmar i ödemarken , så att mitt folk , min utkorade , kan få dricka .
där fanns nämligen en guldsmed , vid namn Demetrius , som förfärdigade Dianatempel av silver och därmed skaffade hantverkarna en ganska stor inkomst .
skapa i mig , Gud , ett rent hjärta , och giv mig på nytt en frimodig ande .
och ännu mycket tydligare blir detta , då nu en präst av annat slag uppstår , lik Melkisedek däri ,
Ty alla de som drivas av Guds Ande , de äro Guds barn .
David själv har ju sagt genom den helige Andes ingivelse : &apos; Herren sade till min herre : sätt dig på min högra sida , till dess jag har lagt dina fiender dig till en fotapall . &apos;
om du framlägger detta för bröderna , så bevisar du dig såsom en god Kristi Jesu tjänare , då du ju hämtar din näring av trons och den goda lärans ord , den läras som du troget har efterföljt .
och vinnläggen eder om att bevara Andens enhet genom fridens band :
därifrån gick den fram österut mot solens uppgång till Gat @-@ Hefer och Et @-@ Kasin och vidare till det Rimmon som sträcker sig till Nea .
då när Gud stod upp till dom , till att frälsa alla ödmjuka på jorden . Sela .
och i vilken man såg profeters och heliga mäns blod , ja , alla de människors blod , som hade blivit slaktade på jorden &quot; .
när han sedan lät Benjamins stam gå fram efter dess släkter , träffade Matris släkt av lotten ; därpå träffades Saul , Kis &apos; son , av lotten , men när de då sökte efter honom , stod han icke att finna .
i veten ju vilka bud vi hava givit eder genom Herren Jesus .
vem mäktar rycka av honom hans pansar ? vem vågar sig in mellan hans käkars par ?
där må prästen Sadok och profeten Natan smörja honom till konung över Israel ; sedan skolen I stöta i basun och ropa : &apos; Leve konung Salomo ! &apos;
och somt föll på stengrund , och när det hade vuxit upp , torkade det bort , eftersom det icke där hade någon fuktighet .
du gör oss till ett trätoämne för våra grannar , och våra fiender bespotta oss .
Nåd vare med eder och frid ifrån Gud , fadern , och Herren Jesus Kristus .
jag skall bliva för Israel såsom dagg , han skall blomstra såsom en lilja , och såsom Libanons skog skall han skjuta rötter .
därför säger HERREN så om konungen i Assyrien : han skall icke komma in i denna stad och icke skjuta någon pil ditin ; han skall icke mot den föra fram någon sköld eller kasta upp någon vall mot den .
Giv mig , min son , ditt hjärta , och låt Mina vägar behaga dina ögon .
Bileam , Beors son , spåmannen , dräptes ock av Israels barn med svärd , jämte andra som då blevo slagna av dem .
därför säger Herren , HERREN Sebaot så : frukta icke , mitt folk , du som bor i Sion , för Assur , när han slår dig med riset och upplyfter sin stav mot dig , såsom man gjorde i Egypten .
när då Husai kom in till Absalom , sade Absalom till honom : &quot; så och så har Ahitofel talat &quot; .Skola vi göra såsom han har sagt ? Varom icke , så tala du &quot; .
hör , dottern mitt folk ropar i fjärran land : &quot; Finnes då icke HERREN i Sion ? är dennes konung icke mer där ? &quot; ja , varför hava de förtörnat mig med sina beläten , med sina främmande avgudar ?
och i din vingård skall du icke göra någon efterskörd , och de avfallna druvorna i din vingård skall du icke plocka upp ; du skall lämna detta kvar åt den fattige och åt främlingen . jag är HERREN , eder Gud .
att man krossar under sina fötter alla fångar i landet ,
i åter skolen icke sluta Förbund med detta lands inbyggare ; I skolen bryta ned deras altaren . &apos; men I haven icke velat höra min röst . vad haven I gjort ! --
den femtonde lotten kom ut för Jeremot , med hans söner och bröder , tillsammans tolv ;
och talen till varandra i psalmer och lovsånger och andliga visor , och sjungen och spelen till Herrens ära i edra hjärtan ,
och när Jehu kom in genom porten , ropade hon : &quot; allt står väl rätt till , du , Simri , som har dräpt din herre ? &quot;
och HERREN har i dag hört dig förklara att du vill vara hans egendomsfolk , såsom han har sagt till dig , och att du vill hålla alla hans bud ;
sedan begav han sig åstad till Tarsus för att uppsöka Saulus .
och Samuel tog sin oljeflaska och göt olja på hans huvud och kysste honom och sade : &quot; se , HERREN har smort dig till furste över sin arvedel .
och Darejaves av Medien mottog riket , när han var sextiotvå år gammal .
hans ben äro pelare av vitaste marmor , som vila på fotstycken av finaste guld . att se honom är såsom att se Libanon ; ståtlig är han såsom en ceder .
Ty deras bördeman är stark ; han skall utföra deras sak mot dig .
och prästerna , leviterna , dörrvaktarna , sångarna , en del av meniga folket samt tempelträlarna , korteligen hela Israel , bosatte sig i sina städer &quot; .
Herren låter höra sitt ord , stor är skaran av kvinnor som båda glädje :
och Josef sade till sina bröder : &quot; jag dör , men Gud skall förvisso se till eder , och föra eder upp från detta land till det land som han med ed har lovat åt Abraham , Isak och Jakob &quot; .
Rikligen mättad är vår själ med de säkras bespottelse , med de högmodigas förakt .
denna sade till sin fru : &quot; Ack att min herre vore hos profeten i Samaria , så skulle denne nog befria honom från hans spetälska ! &quot;
så kan det grönska upp genom vattnets ångor och skjuta grenar lik ett nyplantat träd .
åtta dagar därefter voro hans lärjungar åter därinne , och Tomas var med bland dem . då kom Jesus , medan dörrarna voro stängda , och stod mitt ibland de , och sade : &quot; Frid vare med eder ! &quot;
då skall du svara din son : &quot; vi voro Faraos trälar i Egypten , men med stark hand förde HERREN oss ut ur Egypten .
men en tjänstekvinna , som fick se honom , där han satt vid elden fäste ögonen på honom och sade : &quot; också denne var med honom .
och en man i folkhopen svarade honom : &quot; Mästare , jag har fört till dig min son , som är besatt av en stum ande .
men om en ängel då finnes , som vakar över henne , en medlare , någon enda av de tusen , och denne får lära människan hennes plikt ,
vad man nu därutöver söker hos förvaltare är att en sådan må befinnas vara trogen .
min insikt vill jag hämta vida ifrån , och åt min skapare vill jag skaffa rätt .
Voren I av världen , så älskade ju världen vad henne tillhörde ; men eftersom I icke ären av världen , utan av mig haven blivit utvalda och tagna ut ur världen , därför hatar världen eder .
säg : hör HERRENS ord , du Juda konung , som sitter på Davids tron , hör det du med dina tjänare och ditt folk , I som gån in genom dessa portar .
och han kom till den andre och sade sammalunda . då svarade denne och sade : &apos; ja , herre &apos; ; men han gick icke ,
då sade hon : &quot; se , din svägerska har vänt tillbaka till sitt folk och till sin gud ; vänd ock du tillbaka och följ din svägerska &quot; .
och allt folket och hela Israel insåg då att konungen ingen del hade haft i att Abner , Ners son , hade blivit dödad .
och Jesus sade : &quot; till en dom har jag kommit hit i världen , för att de som icke se skola varda seende , och för att de som se skola varda blinda &quot; .
och detta är lagen om skuldoffret : det är högheligt .
och jag skall föra Israel tillbaka till hans betesmarker , och han skall få gå bet på Karmel och i Basan ; och på Efraims berg och i Gilead skall han få äta sig mätt .
Sjungen till hans ära , lovsägen honom , talen om alla hans under .
eller i det att han , när han har hittat något borttappat , nekar därtill och svär falskt i någon sak , vad det nu må vara , vari en människa kan försynda sig :
av en talent rent guld skall man göra den med alla dessa tillbehör .
de skola sjunga om HERRENS vägar , ty HERRENS ära är stor .
med nardus och saffran , kalmus och kanel och rökelseträd av alla slag , med myrra och aloe och de yppersta kryddor av alla slag .
när bröderna förnummo detta , förde de honom ned till Cesarea och sände honom därifrån vidare till Tarsus .
Foga dem sedan tillhopa med varandra till en enda stav , så att de bliva förenade till ett i din hand .
Jesus svarade och sade till dem : &quot; om jag än vittnar om mig själv , så gäller dock mitt vittnesbörd , ty jag vet varifrån jag har kommit , och vart jag går ; men I veten icke varifrån jag kommer , eller vart jag går .
Käre bröder , bedjen för oss .
men lika lätt kan en dåraktig man få förstånd , som en vildåsnefåle kan födas till människa .
Huru länge , HERRE , skall jag ropa , utan att du hör klaga inför dig över våld , utan att du frälsar ?
då sade han till dem : &quot; från storätaren utgick ätbart , från den grymme kom sötma &quot; . men under tre dagar kunde de icke lösa gåtan .
och om en kvinna i sin mans hus gör ett löfte , eller med ed förbinder sig till återhållsamhet i något stycke ,
Asarja födde Heles , och Heles födde Eleasa .
men Absalom sände ut hemliga budbärare till alla Israels stammar och lät säga : &quot; när I hören basunen ljuda , så sägen : &apos; nu har Absalom blivit konung i Hebron . &apos; &quot;
Herren kom såsom en fiende och fördärvade Israel , han fördärvade alla dess palats , han förstörde dess fästen ; så hopade han över dottern Juda jämmer på jämmer .
ingen som är född i äktenskapsbrott eller blodskam skall komma in i HERRENS församling ; icke ens den som i tionde led är avkomling av en sådan skall komma in i HERRENS församling .
dit Gera jämte Naaman och Ahia förde bort dem : han födde Ussa och Ahihud .
och HERREN sade till Samuel : &quot; Huru länge tänker du sörja över Saul ? jag har ju förkastat honom , ty jag vill icke längre att han skall vara konung över Israel . fyll ditt horn med olja och gå åstad jag vill sända dig till betlehemiten Isai , ty en av hans söner har jag utsett åt mig till konung &quot; .
och alla som bodde i Lydda och i Saron sågo honom ; och de omvände sig till Herren .
de som då togo emot hans ort läto döpa sig ; och så ökades församlingen på den dagen med vid pass tre tusen personer .
åt en gav han fem pund , åt en annan två och åt en tredje ett pund , åt var och en efter hans förmåga , och for utrikes .
när jag alltså vände mig till att jämföra vishet med oförnuft och dårskap -- ty vad kunna de människor göra , som komma efter konungen , annat än detsamma som man redan förut har gjort ? --
och deras barn talade till hälften asdoditiska -- ty judiska kunde de icke tala riktigt -- eller ock något av de andra folkens tungomål .
Ty tre äro de som vittna :
han förde honom fram över landets höjder och lät honom äta av markens gröda ; han lät honom suga honung ur hälleberget och olja ur den hårda klippan .
när de sedan gingo därifrån , bad men dem att de nästa sabbat skulle tala för dem om samma sak .
och han åstundade att få fylla sin buk med de fröskidor som svinen åto ; men ingen gav honom något .
och HERREN gick förbi honom , där han stod , och utropade : &quot; HERREN ! HERREN ! -- en Gud , barmhärtig och nådig , långmodig och stor i mildhet och trofasthet ,
och han sade till honom : &quot; stå upp och gå dina färde . din tro har frälst dig &quot; .
därför har icke heller det förra förbundet blivit invigt utan blod .
och jag , Johannes , var den som hörde och såg detta . och när jag hade hört och sett det , föll jag ned för att tillbedja inför ängelns fötter , hans som visade mig detta .
om däremot allenast få år återstå till jubelåret , så skall han räkna efter detta , sig till godo , och betala lösen för sig efter antalet av sina år .
då sade han till mig : gå ; jag vill sända dig åstad långt bort till hedningarna . &apos; &quot;
och de församlade sig till Jerusalem i tredje månaden av Asas femtonde regeringsår ,
ett mjukt svar stillar vrede , men ett hårt ord kommer harm åstad .
ja , må din hand vara upplyft över dina ovänner , och må alla dina fiender bliva utrotade !
och han sade till dem : &quot; jag har högeligen åstundat att äta detta påskalamm med eder , förrän mitt lidande begynner ;
Ty lika visst som Jesus , såsom vi tro , har dött och har uppstått , lika visst skall ock Gud genom Jesus föra dem som äro avsomnade fram jämte honom .
och när hon har funnit den , kallar hon tillhopa sina väninnor och grannkvinnor och säger : &apos; Glädjens med mig , ty jag har funnit den penning som jag hade tappat bort . &apos;
honom som befaller solen , så går hon icke upp , och som sätter stjärnorna under försegling ;
och alla heliga gåvor som Israels barn giva såsom en gärd , vilken de bära fram till prästen , skola tillhöra denne ;
sedan kallade Abimelek Abraham till sig och sade till honom : &quot; vad har du gjort mot oss ! Vari har jag försyndat mig mot dig , eftersom du har velat komma mig och mitt rike att begå en så stor synd ? på otillbörligt sätt har du handlat mot mig &quot; .
Ty jag vet att I efter min död skolen taga eder till , vad fördärvligt är , och vika av ifrån den väg som jag har bjudit eder gå ; därför skall olycka träffa eder i kommande dagar , när I gören vad ont är i HERRENS ögon , så att I förtörnen honom genom edra händers verk &quot; .
för honom som förvandlar klippan till en vattenrik sjö , hårda stenen till en vattenkälla .
men dessa som stå efter mitt liv och vilja fördärva det , de skola fara ned i jordens djup .
och Jesus begynte åter tala till dem i liknelser och sade :
att de skulle föra drottning Vasti , prydd med kunglig krona , inför konungen , för att han skulle låta folken och furstarna se hennes skönhet , ty hon var fager att skåda .
ja , min boning skall vara hos dem , och jag skall vara deras Gud , och de skola vara mitt folk .
Ty se , de som hava vikit bort ifrån dig skola förgås ; du förgör var och en som trolöst avfaller från dig .
och du skall föra fram hans söner och sätta livklädnader på dem .
och den överskrift som man hade satt upp över honom , för att angiva vad han var anklagad för , hade denna lydelse : &quot; Judarnas konung &quot; .
han skulle ock bliva en fader för omskurna , nämligen för sådana som icke allenast äro omskurna , utan ock vandra i spåren av den tro som vår fader Abraham hade , medan han ännu var oomskuren .
