Om du ansöker om pension från utlandet, får du råd vid Pensionsskyddscentralen.
Kontaktuppgifter till skattebyråns andra serviceställen och telefonrådgivning hittar du på Skatteförvaltningens (verohallinto) webbplats.
Om du vill ha ett arbetsintyg ska du be om det.
Om föräldrarna har ett kombinerat efternamn, blir detta även barnets efternamn.
Skaffa det europeiska sjukvårdskortet i ditt hemland innan du kommer till Finland.
Mer information och råd får du från föreningen Kaapatut Lapset ry.
Att fråga om tillstånd hos hyresvärden om du vill göra ändringar i bostaden, till exempel måla en vägg.
Du får också råd om utarbetandet av en affärsverksamhetsplan och stöd för ditt beslut att starta ett företag.
Om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när hälsostationen öppnar.
Till exempel Sato, Vvo och Avara äger hyresbostäder i Helsingfors.
Oftast betalar hyresvärden förmedlingsarvodet.
Eleverna antas till gymnasiet utifrån vitsorden på avgångsbetyget från grundskolan.
Tolkningfinska
Du kan ansöka till en tionde klass när du har fått ditt avgångsbetyg från grundskolan.
Du kan även registrera bilen på Internet.
Tyvärr kan vi inte svara på respons som är skriven på andra språk.
Företagande kräver yrkeskunnighet och utbildning. Det är viktigt att du är väl insatt i din bransch och lagarna som gäller företagande.
Du kan även besöka mottagningen vid Kliniken för mental- och missbruksvård på servicetorget i Iso Omena utan tidsbokning måndag till fredag kl. 8.30–10.30 och dessutom måndag till torsdag kl. 13–14.30.
Syftet med den partiella sjukdagpenningen är att du kan fortsätta att arbeta eller att återgå till arbetet trots att du har blivit sjuk.
Barnvaktshjälpfinska _ engelska
Du måste beställa tid vid rådgivningarna.
Seure (Seure) är ett bemanningsbolag som erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
Hälsotjänster i Vanda
Om du bor i södra, mellersta eller västra Helsingfors finns hälsocentralsjouren vid Haartmanska sjukhuset.
Ta reda på begränsningarna innan du för in läkemedel i Finland.
Unga i åldern 13–23 med missbruksproblem kan få hjälp vid ungdomsstationen.
personnummer
Kommuninvånarna kan delta i och påverka stadens ärenden vid kommunalvalet som hålls vart fjärde år.
Banken behöver följande uppgifter från dig:
om du ska bo stadigvarande i Finland eller vistas här tillfälligt
Definition av en familj
Giftinformationscentralens telefontjänst är öppen 24 timmar om dygnet.
Med bioavfall avses bl.a.:
Barn vid skilsmässa
Skilsmässa
Den initiala självrisken gäller inte mediciner för personer under 18 år.
krigserfarenheter.
Många organisationer och församlingar bedriver också ungdomsarbete.
Företagsverksamheten startas först när stödet har beviljats.
I Vanda ordnas även många rekryteringsevenemang där arbetsgivarna söker arbetstagare.
Tidsbokningen kan du ringa:
Anmälan utan nätbankskoderfinska _ svenska
Lapplands universitetfinska _ engelska
Gymnasiestudierna siktar till studentexamen (ylioppilastutkinto).
Varken staden eller andra hyresvärdar har skyldighet att erbjuda dig bostad.
Vid hälsostationernas preventivrådgivning (ehkäisyneuvola) får du hjälp med graviditetsprevention och familjeplanering.
Din chef berättar för dig om du behöver ett läkarintyg om sjukdomen direkt eller först från och med den fjärde sjukledighetsdagen.
Våld Problem i äktenskap eller parförhållande
Flerspråkiga biblioteketfinska _ svenska _ engelska
bilda ett kombinerat efternamn av era efternamn.
du är medborgare i ett EU-land, EES-land eller Schweiz och du har
Du kan få kostnadsfri hjälp vid Kyrkans familjerådgivningscentral även på engelska och svenska, även om du inte är medlem i kyrkan.
Teatrar i Esbofinska _ svenska _ engelska
På utbildningsstyrelsens (opetushallitus) webbplats finns en sökmotor med vilken du kan se var och när du kan avlägga examen.
Även minderåriga barn kan boka tid hos läkaren och få ett recept för preventivmedel.
Spara lönekvittona.
Mer information om sport som hobby hittar du på InfoFinlands sida Motion.
linkkiMarthaförbundet:
Tandvårdens tidsbeställning och värkjouren nås vardagar kl. 8–15 på tfn 016 322 2562 eller 016 356 1750. Kvällstid och på veckoslut kan du ta kontakt med läkarmottagningen om du är i brådskande behov av vård.
Vid Grankulla konstskola kan barn och unga studera bildkonst och vid Grankulla musikinstitut kan barn och vuxna studera musik.
Min arbetsgivare hotar mig dessutom med våld.
Äldre människors hälsa, Äldre människor
I Finland anlitar många företag revisionsbyråer.
Partiell förtida ålderspension
Mer information om ledigheterna får du på InfoFinlands sida Familjeledighet.
som en kyrklig vigsel.
Erkännande av examen är avgiftsbelagt.
Processen är mycket snabb och smidig.
Om du bor i höghus eller radhus ska du alltid också komma ihåg att meddela husets disponent (isännöitsijä) att du flyttar.
En demonstration ska anmälas till polisen på förhand.
linkkiFörbundet Utvecklingsstörning:
Fundera noga hur företaget drivs och var och hurdana lokaler företaget har.
Seniorrådgivningenfinska _ svenska
Flyktingstatus får de som beviljas asyl eller som tas till Finland i flyktingkvoten.
Kommunerna
Jobben finns till exempel på skolor, daghem och sjukhus.
Arbete med ett annat uppehållstillstånd
bor permanent i Finland
du är arbetslös eller kommer att bli arbetslös
Tolken ska vara vuxen, egna minderåriga barn kan alltså inte användas som tolk.
Könssjukdomar behandlas i huvudstadsregionen på polikliniken för könssjukdomar i Helsingfors.
Karleby evangelisk-lutherska församlingar erbjuder även hobbyverksamhet för barn och unga, såsom lekparksträffar, klubbar, musikverksamhet och läger.
Avgiftens storlek beror på hur många böcker som är försenade och hur många dagar de är försenade.
Också företagaren har rätt till utkomstskydd för arbetslösa.
Därefter placeras invandrareleverna i en finskspråkig klass i sin närskola.
Du kan också bo hemma och gå på rehabilitering därifrån.
Kandidaten ska vara en person
Om du behöver information om hälsotjänsterna, kan du ringa hälsorådgivningen: (09) 310 100 23.
Vistelsetiden på tre månader räknas alltid från det att du varit utanför Finlands gränser.
Möjligheter att studera det finska eller svenska språket
Arbetarskyddsmyndigheten kan förplikta arbetsgivaren att rätta till brister i arbetssäkerheten som förekommer på arbetsplatsen
Lägg till kontaktuppgifterna till dem.
Förskoleundervisning
Kontakta magistraten på din hemort om meddelandet om rösträtt inte skickas hem till dig.
Observera att listan inte nödvändigtvis innehåller allt som måste göras när du flyttar till Finland.
Fpa:s stöd för boendet är följande:
Som fristående examen (näyttötutkinto) (vuxenstuderande)
Arealen är cirka 240 km2, varav cirka 2 km2 består av vatten.
Gymnasieskolorfinska
Kommunerna tillhandahåller många tjänster för sina invånare.
Enligt lag får man inte beställa läkemedel per post från länder utanför EES-området.
Vid problem hos unga i skolåldern hjälper exempelvis skolans hälsovårdare eller skolkuratorn.
Du får hjälp med jobbsökningen på arbets- och näringsbyrån (Työ- ja elinkeinotoimisto), d.v.s. TE-byrån.
Delta och påverkafinska _ svenska _ engelska
Föreningar och organisationer samt hobbygrupper och kommunala institut erbjuder kurser i idrott och kultur samt bl.a. språk och hantverk.
Om du själv bokar tolken och betalar kostnaderna kan du anlita en tolk när som helst.
Skriv ut blanketten på Migrationsverkets webbplats och fyll i den färdigt.
dina rättigheter och skyldigheter
Vem som helst kan ansöka om ett bostadslån hos banken.
Ekonomi- och skuldrådgivningfinska.
I InfoFinland under rubriken Officiellt intyg över språkkunskaper får du information om hur du kan jämföra kursernas nivåer med nivån på den allmänna språkexamen (yleinen kielitutkinto).
Examen vid sidan av arbetet med läroavtal
Verksamhetsställen för handikappservicefinska
Du behöver ändå inte borgensmän för ditt lån om du har sparat ihop en del av bostadens pris på förhand, eller om du har annan egendom som duger som säkerhet för lånet.
Läs mer: När du väntar barn.
Klamydia och gonorré behandlas med antibiotika.
Om du inte är kund hos en mottagningscentral kan du ansöka om stöd hos Migrationsverket.
I de lägre årskurserna har man cirka 20 undervisningstimmar i veckan och antalet ökar i de högre årskurserna.
Dessutom har vissa läroanstalter egna studenthem.
Medborgarinstitut
Information för utländska studerandeengelska
legitimation (till exempel pass)
Öppen ansökan
Hälsovårdscentralen
Du får mer information om rätten till hemkommun på InfoFinlands sida Hemkommun i Finland.
Medier
barn och föräldrar
Teater
ortodoxa kyrkan (ortodoksinen kirkko) eller
Därför skulle det vara bra att barnen hade möjlighet att röra på sig tillräckligt också utanför daghemmet eller skoltiden.
Lagar och avtal i arbetslivet
En utredning om dina språkkunskaper
linkkiJämställdhetsombudsman:
På hälsostationen behandlas de vanligaste psykiska problemen.
KOSEK (Karlebynejdens Utveckling Ab) erbjuder tjänster som nyttar företaget under hela dess livscykel, från och med att starta företagsverksamhet.
I Vanda finns också många andra hyresvärdar, varav de största är VVO, Sato och Avara.
Man kan inte heller föreslå en annan person, till exempel en släkting eller vän, som kvotflykting.
Samtal till huvudhälsostationen styrs till ett och samma telefonnummer, (06) 8287 310.
Adress: Steniusvägen 20, 00320 Helsingfors
de som bor i kollektiv.
Transsexuella personer, transvestiter, intersexuella personer och andra människor med mångfacetterad könsidentitet kan få hjälp av jämställdhetsombudsmannen om de upplever diskriminering.
Stadin ammattiopisto är Finlands största yrkesläroanstalt där man kan utbilda sig inom många olika branscher.
Flyttjänsterfinska _ engelska _ ryska
Hälsostationerna har öppet måndag till fredag kl. 8–16.
Information om anmärkning om betalningsstörningfinska _ svenska _ engelska
Handikappservice och stödåtgärderfinska _ svenska _ engelska
Huruvida du omfattas du av den sociala tryggheten och kan få bidrag påverkas också av om du flyttar till Finland till exempel som
Guiden Välkommen till Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska
Om du orsakar skador i bostaden måste du ersätta dem.
Läs mer på InfoFinlands sida Yrkesutbildning.
På stadens webbplats finns information om stadsfullmäktige och dess beslut.
Vård av barn i hemmetfinska _ svenska _ engelska
Information om konsumenträttigheterfinska
yrkesvägledning
Om du söker arbete, bör du anmäla dig till TE-byrån.
Du får närmare uppgifter vid social- och närarbetets verksamhetsställe i ditt bostadsområde (sosiaali- ja lähityön toimipiste).
Appar
Grundskolans övriga stödåtgärder omfattar den övriga stödundervisningen i grundskolan, specialundervisning, individuella studieplaner, flexibel bedömning,
Var kan jag få hjälp?
Information om riksdagenfinska _ svenska _ engelska
Om du är under 16 år och behöver preventivmedel, ta kontakt med hälsovårdaren vid din läroinrättning.
Du får personbeteckningen, när du registrerar dig som invånare hos magistraten.
Diskrimineringsombudsmannens kundtjänstfinska _ svenska _ engelska
Om du har ett tillfälligt uppehållstillstånd (B-tillstånd) som är i kraft kan du få en hemkommun om du kan påvisa att det är din avsikt att bo stadigvarande i Finland.
I lågstadiets högre klasser och på högstadiet får de även välja tillvalsämnen.
Inrikesministeriet beslutar från vilka länder kvotflyktingarna tas.
Om samborna har gemensamma minderåriga barn ska de tillsammans besluta om barnens situation på samma sätt som vid skilsmässa.
Många saker i det finländska samhället förändrades.
Om du inte är säker på huruvida banken ger dig ett lån lönar det sig att gå till banken och förhandla om lånet i god tid innan du köper bostaden.
Du ansöker om visum med en visumansökningsblankett.
I samma lokal finns kundtjänsten Osviitta, där du kan köpa resekort till lokaltrafiken.
I vissa gymnasier ges även mycket undervisning i konstämnen.
Från länder utanför EES-området får du ta med dig till Finland den mängd läkemedel för eget bruk som motsvarar högst tre månaders förbrukning.
Navigatorns Startpunkter erbjuder handledning och rådgivning utan tidsbokning till unga under 30 år.
Webbplatsen asuminen.fifinska _ svenska _ engelska
Studentbostäder hyrs ut av studentbostadsstiftelser, universitetens studentkårer, nationer och vissa andra stiftelser.
Du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv.
Klockan 8.00 betyder prick klockan 8.00, inte klockan 8.10.
Vem kan rösta?
Om du brådskande behöver hjälp av Polisen i en nödsituation ska du ringa nödnumret 112.
Enligt Finlands lag är män och kvinnor jämställda.
Du kan göra en anmälan om medborgarskap på internet.
Norrskenfinska _ engelska
Vid skilsmässa kommer man överens om hos vilken förälder barnet har sin officiella adress.
Undervisning i det egna modersmålet för invandrare
Skatteförvaltningen gör en del avdrag automatiskt, men vissa avdrag måste du själv ansöka om.
Om du har det europeiska sjukvårdskortet (European Health Insurance Card, EHIC), behöver du ingen separat försäkring.
Sök till högre yrkeshögskolestudier i den gemensamma ansökan.
Allmänt om fackförbund
Du kan få rehabilitering om ditt handikapp orsakar stora svårigheter att klara av vardagen i hemmet, skolan eller arbetet.
En annan anhörig kan få uppehållstillstånd också om han eller hon levt tillsammans som en familjemedlem till den anhöriga som är bosatt i Finland, innan denna person kom till Finland.
Utbildning för invandrarefinska
Lapplands arbets- och näringsbyrå
Vatten
Till slut anslöts hela Finland år 1809 till Ryssland, efter att Ryssland besegrat Sverige i krig.
Mer information om reglerna i Finland ges av Livsmedelsverket (Ruokavirasto).
Läs mer: Brott.
Läs mer om att grunda ett företag på InfoFinlands sida Att grunda ett företag.
Utbetalningen av semesterpenning baserar sig på kollektivavtalet.
du startar företagsverksamheten först när stödet har beviljats.
För ett bostadslån behövs det vanligen en säkerhet (vakuus).
68300 Kelviå
Ofta kan du utbilda dig på arbetstid och arbetsgivaren kan betala för utbildningen.
vård för att förbättra arbets- och funktionsförmågan
Du kan också göra ditt slutarbete i något företag eller göra en arbetspraktik.
Hjälptelefon: 020 316 116
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
När du ansöker om det första uppehållstillståndet i Finland kan du även be om registrering i det finska befolkningsdatasystemet.
Synskadade
Läs mer på InfoFinlands sida Finska och svenska språket.
Skatteprocenträknarefinska _ svenska _ engelska
Tidpunkten varierar men oftast firas påsk i mars eller april.
Morsdag
Via Wilma kan du ha kontakt med barnets lärare och få information om barnets lärande, prov och frånvaron samt händelser i skolan och om skollov.
Sök en bostad i god tid innan du flyttar till Finland
Arbetsgivaren kan även betala handläggningsavgiften för arbetstagaren.
Barnet får automatiskt finskt medborgarskap vid födseln i följande fall:
I detta fall ska du ansöka om en finsk personbeteckning och meddela din adress till magistraten (maistraatti).
Mer information om personbeteckningen hittar du på InfoFinlands sida Registrering som invånare.
Aktiebolaget är den vanligaste företagsformen i Finland.
Bröstcancerundersökningen görs för kvinnor i åldern 50–69 år ungefär vartannat år och undersökningen för livmoderhalscancer för kvinnor i åldern 30–60 år med fem års mellanrum.
Kontrollera vilket alternativ som är förmånligast för dig.
Med hjälp av tjänsten finnishcourses.fi kan du söka en lämplig kurs i finska i Helsingfors, Vanda, Esbo eller Grankulla.
I detta fall måste du göra en underrättelse om rörlighet till Migrationsverket.
Bland annat hos bostadsförmedlingen, på internet och i lokala tidningar finns annonser om bostäder som är till salu.
Utländska medborgare
Finlands kulturhistoria kan du bekanta dig med bland annat i Finlands nationalmuseum som ligger i Helsingfors.
Läs mer: Teater och film.
Den kostnadsfria rådgivningen ges på finska och engelska.
Ungdomar kan diskutera frågor kring sexuell hälsa med hälsovårdaren vid sin egen skola.
I Helsingfors finns gott om cykelvägar.
Ubildning vid öppna universitetet i Vandafinska _ svenska _ engelska
På Navigatorn kan någon i personalen hjälpa dig att reda ut saker och ting.
Lägenhetshyrorna är vanligen i genomsnitt 100 euro per dygn.
Därtill utbetalas barnbidrag (lapsilisä) till barnets vårdnadshavare fram till dess att barnet fyller 17 år.
Du hittar anvisningar och mer information om ansökan om uppehållstillstånd för uppstartsföretagare på Migrationsverkets och Business Finlands webbplatser.
Asylsamtalet (turvapaikkapuhuttelu) är den viktigaste händelsen under behandlingen av din ansökan.
Till exempel befinner sig en studerande vars enda orsak till vistelsen i landet är studierna tillfälligt i Finland.
Kommunernas idrottsplatser får användas av alla invånare.
På InfoFinlands sida Var hittar jag jobb? finns information om hur du kan hitta ett jobb i Finland.
Dessutom kan du få stöd, rådgivning och handledning.
Läs mer på InfoFinlands sida Barns och ungas problem.
Karlebynejdens institut, som ägs och drivs av Karleby stad, är ett tvåspråkigt (finska och svenska) medborgarinstitut.
Egenvårdsläkemedel (itsehoitolääke) kan köpas utan läkarrecept.
Mer information om makarnas egendom hittar du på InfoFinlands sida Äkta makars rättigheter och skyldigheter.
Rådgivning för och integration av invandrare
Läs mer på InfoFinlands sida Barn vid skilsmässa.
Arbetsgivaren utser för varje arbetsplats en arbetarskyddschef, som bistår arbetsgivaren i samarbetet med anställda och arbetarskyddsmyndigheter.
Om du har anställning i Finland, är det skäl för dig att ansluta dig till en finländsk arbetslöshetskassa.
Om du är studerande kan du söka hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS.
Bibliotekstjänsterfinska _ svenska _ engelska
Läs mer: Yrkeshögskolor, Universitet.
nivåerna B1 och B2: en självständig språkanvändares språkkunskaper (itsenäisen kielenkäyttäjän kielitaito)
Du får då avdragen i efterskott som en skatteåterbäring.
Medlemskapet i panelen binder dig inte till någonting.
Målet är att främja hälsan och välbefinnandet för de blivande föräldrarna och hela familjen och att stöda familjen inför deras nya uppgift som föräldrar och i växelverkan.
Video om arbetstagarens rättigheter i Finlandengelska _ kinesiska _ arabiska _ thai _ hindi
Hyresbostad
Avfallsinsamlingsstationerfinska
På InfoFinlands sida Val och röstning i Finland finns information om vem som kan rösta i kommunaval.
På arbetsplatser och i skolor serveras lunch vanligtvis kl. 11–12.
Vem som helst kan behöva hjälp om livssituationen är påfrestande.
De är fel som ingen känner till.
Centraliserad tidsbokning per telefon: (06) 8287 400
Församlingarfinska _ svenska
Uppsägning av hyresavtal
Se till att det finns tillräckligt många brandvarnare i ditt hem.
Det är bra att skaffa sig en Internetuppkoppling så fort som möjligt efter att du har flyttat till Finland.
På denna sida finns information riktad till kvotflyktingar.
I Helsingfors kan du bli kund hos rådgivningen om du har ett FPA-kort.
Detta innebär att de inte har rätt till FPA:s förmåner.
Fråga mer vid din förläggning.
Du kan också avsluta studierna efter lägre högskoleexamen.
finns information om hur du kan hitta ett jobb i Finland.
Evenemang i Grankullafinska _ svenska _ engelska
Om din hemkommun är Vanda kan du använda kommunens offentliga hälsovårdstjänster.
skattekort och skattenummer samt rådgivning om beskattningen
Om du arbetar vid sidan av studierna är din arbetstid begränsad.
Spara intygen från dina tidigare jobb och studier.
Dessa dagar kan du dela upp på högst fyra perioder.
Läraren bedömer elevernas framsteg i skolan.
Allmän språkexamen, ASE, är ett språktest för vuxna.
Barn som har ett annat modersmål än finska eller svenska kan få modersmålsundervisning.
Vanda erbjuder ungdomar under 20 år gratis preventivmedel.
Webbaserat material
Dagvård i Helsingforsfinska _ svenska _ engelska
Lapplands yrkesinstitut
Trafikfinska _ svenska _ engelska
Information om Migrationsverketfinska _ svenska _ engelska
På finska duar man oftast.
Det är viktigt att du beskriver allt som hänt så exakt som möjligt.
Många städer har rådgivningstjänster för invandrare med rådgivare som specialiserat sig på invandringsfrågor.
Om du bor i en hyresbostad ska du komma ihåg att säga upp din gamla bostad i tid.
Rysktalande klienter: 020 634 4901 (mån.–fre. kl. 10–12 och 13–15)
Läs mer: Trafik.
Det är bra om paret besöker mottagningen tillsammans.
minst tre års arbetserfarenhet från en lämplig bransch
Om man vill fortsätta studierna därefter och avlägga högre yrkeshögskoleexamen, måste man först skaffa sig tre år av arbetserfarenhet från samma område som examen.
Jag måste flytta ut på grund av skilsmässa.
Information om gymnasiestudierfinska _ svenska
De viktigaste verksamhetsformerna består av ungdomsgårdarna, stora ungdomsevenemang, utflykter, internationella utbyten för ungdomsgrupper och sommarkollon för barn.
kursanmälanfinska
Områdeskoordinatorn berättar om hur undervisningen ordnas och hjälper dig i frågor som rör barnets skolgång.
Bostadsrättsbostäderfinska _ svenska _ engelska
Finland för att bo hos en familjemedlem ska du ansöka om registrering av uppehållsrätten för EU-medborgare på grund av familjeband i tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Befolkning
Åldringar
På magistraten utreder man om det är möjligt att registrera en hemkommun (kotikunta)för dig.
Du har rätt att använda arbets- och näringsbyråns tjänster om du har fått kontinuerligt uppehållstillstånd (A) eller permanent uppehållstillstånd (P).
Du kan dra av låneräntan i beskattningen.
Om arbetsavtalet är tidsbundet binder det båda parterna en bestämd tid, om man inte har kommit överens om möjligheten till uppsägning.
På webbplatsen för MIELI Psykisk Hälsa Finland rf (MIELI Suomen Mielenterveys ry) hittar du information om
festivalarbete
Barnet kan även delta i småbarnspedagogik tillsammans med föräldern i lekparker.
P-EU-tillståndsansökan kan även avslås på samma grunder som permanent uppehållstillstånd.
Du behöver följande handlingar:
Videoklipp och broschyrer för invandrarefinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska
LaNuti linkkiLaNuti:
Information om boendefinska _ engelska
Då är tolkningen kostnadsfri för dig.
Skilsmässa och vårdnad om barn
Överväger du att avbryta graviditeten?
Du krävs inte på redogörelse över din utkomst.
linkkiCIMO:
Läs mer: Stöd- och serviceboende
Det finns också caféer där kunderna har möjlighet att använda Internet.
Nationalparkerfinska _ svenska _ engelska _ ryska _ kinesiska
sexuell läggning.
I början av CV:t kan du tillfoga en sammanfattning eller profil där du beskriver din bakgrund och din kärnkompetens med några ord.
Finskans grammatikengelska
På den här sidan finns information om tjänsterna i Rovaniemi.
Chatbot-tjänst för utländska företagarefinska _ engelska
Påsk
Bästa stället att fråga om enskilda grenar och var man kan utöva dem är grenförbunden.
Ta med dig identitetsbevis och uppehållstillstånd.
Sporrgränden 2 A, vån. 3 (Håkansböle)
Du kan också vända dig till Huvudstadens Skyddshem (Pääkaupungin Turvakoti).
FPA ordnar rehabiliteringen och ersätter kostnaderna för den.
Privat psykoterapitjänst på Internetfinska _ svenska _ engelska _ ryska _ franska _ spanska _ turkiska _ kinesiska _ tyska _ portugisiska _ norska
En brandvarnare kan rädda ditt liv.
Barn kan också gå i en skola med en speciell inriktning.
Hen ger dig råd och ser till att dina rättigheter förverkligas.
När en person som är fast bosatt i Finland blir arbetslös, har han eller hon rätt att få utkomstskydd för arbetslösa.
Förmånligast övernattar man i delat rum.
Bostäderna är dyrare nära stadens centrum.
Om man bryter mot trafikreglerna kan man få böter.
Finland accepterade resedokumentfinska _ svenska _ engelska
Arbetsgivaren kan ansöka om stöd för arbetstagarnas finskundervisning via arbets- och näringslivstjänsterna.
Skyddshemmet Mona är endast avsett för invandrarkvinnor och deras barn.
De offentliga tjänsterna började utvecklas och på så sätt skapade man den offentliga hälsovården, sociala tryggheten och grundskolan.
För att kunna ansöka om ett nytt uppehållstillstånd för arbetstagare måste du ha ett nytt jobb.
Kindpussar är dock ovanliga.
Dixi, Banvägen 11, 2:a vån.
Du kan prata om dina problem med skolans eller läroanstaltens hälsovårdare eller de vuxna vid ungdomsgården.
Om du vill kan du även be någon annan släkting eller en vän att följa med.
En utvecklingsstörd person som behöver vård kan bo i ett familjehem.
Lapplands yrkesinstitut
tfn (09) 8392 3415
På universitet kan man avlägga lägre högskoleexamen på cirka tre år och därefter högre högskoleexamen på cirka två år.
Helsingfors stad ordnar eftermiddagsverksamhet för barn i årskurs 1 och 2 i skolor och lekparker efter skoldagen.
Tfn 029 55 39391
Myndigheterna överväger beviljandet av uppehållstillstånd alltid fall för fall.
Detta kallas för aktiveringsmodellen för arbetslöshetsförsäkringen (työttömyysturvan aktiivimalli).
Du får stanna i Finland om du beviljas asyl eller uppehållstillstånd på någon annan grund.
Du kan lära dig ett nytt yrke eller en ny examensdel.
Regler
Ansvarig bolagsman i kommanditbolag
Finlands utrikespolitik i samverkan med statsrådet och
Grundläggande information om yrkeshögskolorfinska _ svenska
Du har möjlighet att få en hemkommun i Finland om:
Dessa nivåer delas ytterligare in i undernivåer.
Passfoto (anvisningar för fotot finns på Migrationsverkets webbplats)
På hjälptelefonen får du stöd och vid behov råd om var du kan få hjälp.
Konserterfinska _ svenska _ engelska
Privata mentalvårdstjänster
Läs mer: Högskoleutbildning.
Företagsverksamhet som bisyssla lönar det sig ofta att starta som enskild näringsidkare.
Separat insamlat bioavfall packas i en papperspåse, en påse vikt av en dagstidning eller en plastkasse. Kassen eller påsen får vara högst 30l stor.
Invånarhusen Kivenkolo och Kylämaja är öppna för alla.
För dessa koder gäller dock hårdare krav än för öppning av ett bankkonto.
Du kan även söka fram en privat advokat via Finlands Juristförbunds webbplats.
Om bostaden är större eller dyrare än vad lagen om allmänt bostadsbidrag tillåter växer den andel av boendekostnaderna som du betalar själv.
För att teckna ett abonnemang behöver du ett finländskt identitetsnummer och du måste ha en adress i Finland.
På utbildningsstyrelsens (opetushallitus) webbplats finns en sökmotor för språkexamina.
Öppet varje dag dygnet runt.
Bildkonst
Dessutom krävs att:
Ta i god tid reda på när du kan ansöka om en studieplats.
Övriga länders medborgare måste anmäla sig personligen hos TE-byrån.
Då ordnas fyrverkerier.
Kvinnan har rätt att själv besluta om hon vill göra abort.
Då kan domstolen döma till skilsmässa direkt.
Hur ordnas umgänget?
En besvärsanvisning om hur beslutet får överklagas bifogas alltid beslutet.
Läs mer om sjukförsäkringen i Finland på InfoFinlands sida Den sociala tryggheten i Finland.
Utbudet kompletteras av språk- och metodstudier.
I hälsovården av barn under skolåldern får man hjälp av rådgivningsbyråerna (neuvola).
Diskriminering (syrjintä) är ett brott.
På Finlex webbplats kan du läsa lagen angående vårdnad om barn och umgängesrätt.
Studierna omfattar mycket praktiska övningar.
Privat dagvårdfinska
Telefon: 029 56 49294
Vid vårt vetenskaps- och konstuniversitet fås utbildning och idkas forskning inom pedagogik, turism och affärsverksamhet, juridik, konstindustri och samhällsvetenskaper.
Europass är särskilt nyttigt om du ansöker om ett jobb eller en utbildningsplats i Finland från ett annat EU-land.
När du ansluter dig till ett fackförbund kan du samtidigt ansluta dig till förbundets arbetslöshetskassa.
Det finns inga möjligheter att övernatta på nattcaféet, och det är inte heller drogfritt.
Hälsostationernas adresser:
Du kan använda de offentliga hälsovårdstjänsterna om du har en hemkommun i Finland.
På InfoFinlands sida Att grunda ett företag hittar du information om hur man grundar ett företag i Finland.
För hormonella preventivmedel behöver du ett recept av en läkare.
Familjeledigheter
Hälsostationen på Rinteenkulmafinska
Också sökandens inkomster beaktas, eftersom bostäderna främst är avsedda för personer med låga inkomster.
Utbildning som handleder för yrkesutbildning (VALMA)
Samhället tryggar barnets rättigheter med hjälp av lagar och författningar.
Enligt Finlands lag ska alla människor behandlas likvärdigt oberoende av deras bakgrund och kön.
Det åligger kommunerna att ordna serviceboende och stödboende för personer som behöver det.
Du kan ta direkt kontakt med en arbetsplats som du är intresserad av.
Läs mer:
Ibland är dessa skolor privatskolor.
Finska medborgares rättigheter och skyldigheterfinska _ svenska _ engelska
Din uppehållsrätt kan registreras om du är anställd eller har ett eget företag i Finland.
Det har på grund av förälderns ekonomiska situation fastställts att inget underhållsbidrag betalas.
Avtala om arvodet skriftligen på förhand.
Studentexamen består av prov i olika läroämnen.
Du får alltså både yrkesutbildning och en arbetsplats.
Juristens rådgivning per telefon 020 316 117
Diabetes kan behandlas med insulin och rätt kost.
Att röra sig i naturen
Förete skattekortet till din arbetsgivare.
Mer information hittar du på FPA:s webbplats.
Hyresbostäderfinska _ svenska
hör till en finländsk arbetslöshetskassa
Vid Esbo musikinstitut (Espoon musiikkiopisto) kan barn och vuxna studera musik.
du har tidigare haft en hemkommun i Finland
I staden finns flera busslinjer.
De flesta utrikesflygen avgår från Helsingfors-Vanda flygplats.
Läs mer på InfoFinlands sida Dödsfall.
Kasta inte avfallet ut genom fönstret, i skogen eller på gatan.
Du hittar jobbförmedlingssidor när du skriver "avoimet työpaikat" (lediga jobb) i sökmotorns sökfält.
Migrationsverket skickar dig en kallelse till asylsamtal.
De högsta tjänstemännen i Rovaniemi stad är stadsdirektören och två biträdande stadsdirektörer.
I Finland kan du studera på finska, svenska och ibland på engelska.
Sådana preventivmedel är till exempel p-piller och minipiller.
Förskoleundervisningen är avsedd för sexåringar och den ges vid daghem.
När du har en hemkommun kan du använda kommunens tjänster, såsom till exempel hälsovårdstjänster.
ryska och engelska tfn 050 325 7173
Det allmänna nödnumret är 112.
Om du är sambo med en finsk medborgare som bor i Finland kan du få uppehållstillstånd på grund av familjeband.
Du kan även ta dig till Huvudstadens Skyddshem.
Evenemang och sevärt i Helsingforsfinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Söka bostad
Ainonkatu 1, vån.
Enligt lag får ingen diskrimineras till exempel av följande orsaker:
Att ansöka om skilsmässa
Du får mer information om tolktjänsterna i din kommun på rådgivningsbyrån.
Presidentval
Låt göra en läkarundersökning före utgången av den fjärde graviditetsmånaden.
När Migrationsverket har gett ett positivt beslut på din ansökan om återförening på grund av familjeband och anser att staten kan bekosta resan för dina familjemedlemmar, skickar det sitt beslut till Röda Korset.
Observera att tull- och skattefriheten för flyttsaker inte gäller alkohol eller tobaksprodukter.
Motion
Till reglerade yrken hör både uppdrag inom den offentliga sektorn och yrken för vilka det krävs rätt till yrkesutövning.
Du kan studera finska eller svenska.
Då firas i Finland midsommar, som är midnattssolens och högsommarens fest.
En utredning om ditt uppehälle.
På Omnia ordnas för invandrare utbildning som förbereder dem på yrkesutbildning.
Nylands arbets- och näringsbyrå, Esbo
vistas i landet illegalt
I arbetslivet ska kvinnor och män behandlas lika.
Tfn (09) 839 21074 och (09) 839 32042
Vuxna invandrare som inte har grundskolans avgångsbetyg från sitt eget land kan avlägga grundskolan på vuxengymnasiet.
Det kan variera allt mellan dagliga till veckovisa hembesök.
Nollalinja är en hjälptelefon som du kan ringa om du har blivit utsatt för våld i familjen, sexuellt våld eller hot om våld.
Barnskyddslagen (Lastensuojelulaki) säger att alla barn bosatta i Finland har rätt till omsorg och en trygg uppväxtmiljö.
Rehabiliterande psykoterapifinska _ svenska _ engelska
Företagare som säljer varor och tjänster i Finland är skyldiga att betala mervärdesskatt.
Fångstvägen 3
Bio Rex program finns under länken här intill.
Vid yrkeshögskolorna och universiteten i Esbo och Helsingfors kan du studera inom många områden.
rehabiliteringspsykoterapi
Om du blir arbetslös
Studierna på studielinjerna pågår i 1–2 år.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kontakta ett skyddshem.
Människohandelns offer kan få hjälp.
Om du inte korrigerar skattedeklarationen, förblir det här beskattningsbeslutet i kraft.
Om du inte betalar räkningen senast på förfallodagen eller inte har kommit överens om att förlänga betalningstiden, måste du betala påminnelse- och inkassokostnader samt dröjsmålsränta.
Exporten av tjära, som blev mycket viktig för Karlebys historia, inleddes redan på 1500-talet.
Att köpa sexuella tjänster av ett barn under 18 år är ett brott.
Tidsbeställning
Största delen av läkemedelsbutikerna på internet är dock illegala.
Om du har en funktionsnedsättning, ta då först kontakt med hälsostationen (terveysasema).
Velkalinja är Takuusäätiös kostnadsfria rådgivningstelefon.
67701 Karleby
Meddela numret på ditt bankkonto via Skatteförvaltningens webbtjänst eller på en separat pappersblankett.
Intern kommunikation på arbetsplatsen
Av det ser arbetsgivaren, hur mycket skatt som ska betalas på lönen.
Den är gratis.
Finlands förhistoria –1323
På InfoFinlands sida Våld hittar du information om vad du kan göra om din partner utövar våld eller hotar med våld.
Du måste meddela daghemmet och skolan när barnen slutar där.
Mariegatan 16–20 (l-flygeln, ingång B1)
Hyresvärden har hotat med att vräka mig från hyresbostaden på grund av högljutt liv.
Kvällar och helger
Du kan söka till en yrkesutbildning när du har avlagt lärokursen för den grundläggande utbildningen.
Etableringsanmälan
Läs mer: Hyresbostad.
Om din närstående utgör en fara för sig själv eller för andra och inte går med på att träffa en läkare kan du ringa hälstocentralen eller sjukhuset.
Förlossningfinska _ svenska _ engelska
Polikliniken för könssjukdomarfinska _ svenska _ engelska
Om säljaren av bostaden godtar köpeanbudet görs bostadsköpet upp i köparens bank.
Mer information om möjligheter till musikhobby får du via kommunens kulturkontor.
Den internationella föreningen i Håkansböle (Hakunilan kansainvälinen yhdistys) har en rådgivningspunkt som betjänar invandrare i Håkansböle, Björkby och andra områden i Vanda, som vill ha information om till exempel studier, språkkurser, arbete, hobbyverksamhet, krissituationer eller juridiska frågor.
Du kan inte få flexibel eller partiell vårdpenning om du får föräldradagpenning och/eller hemvårdsstöd och själv tar hand om dina barn.
Folket kom österifrån från nuvarande Rysslands område och söderifrån via Baltikum.
Karleby finska gymnasium erbjuder förberedande undervisning för gymnasiet även för invandrare.
omfattas av den finländska sjukförsäkringen (sairausvakuutus): läs mer på InfoFinlands sida Den sociala tryggheten i Finland
Information om finska romanifinska
På daghemmet är barnen i större gruppen är i gruppfamiljedagvården.
Folk flyttar till Finland
Delägare som innehar en ledande ställning i ett aktiebolag (verkställande direktör eller styrelsemedlem) eller person som innehar en ledande ställning i någon annan sammanslutning
Skrapning görs vanligtvis i narkos och därefter ska du stanna några timmar på sjukhuset.
Måste jag betala?
Du kan även fråga om mer information av daghemsföreståndarna.
Minnesstörningar och demensfinska _ svenska _ engelska
Fråga om råd på företagsrådgivningen
dina inkomster inte är för stora; och
FPA
Den närmaste byrån finns i Esbo.
Man kan ansöka om bodelningsman om samboförhållandet har varat minst fem år och parterna har gemensamma barn.
Gymnasiet är en allmänbildande utbildning som inte ger ett yrke.
Publikationer eller andra arbetsprov
Tfn 09 3104 4556 (mån–fre kl. 9–15)
Familjerådgivningscentralenfinska
På stadens webbplats hittar du också anvisningar om hur du söker hyresbostad.
Finskt medborgarskap till barn med finsk farfinska _ svenska _ engelska
Bostadsrättsbostäderfinska
linkkiMetropolia:
Finnkino är den största biografkedjan i Finland.
När du blir sjuk ska du kontakta hälsostationen i ditt område.
Barnkulturcentralen Musikantitfinska _ engelska _ ryska
En studerande från ett land utanför EU/EES kan ha rätt till vissa av FPA:s förmåner, till exempel de förmåner som ingår i sjukförsäkringen.
Hörselapparatfinska
Läs mer: Hälsovårdstjänster i Finland.
Stöd för familjer
Om du utsätts för diskriminering kan du be om hjälp av Diskrimineringsombudsmannen.
Hälsa och rehabiliteringfinska _ svenska _ ryska _ estniska
De ungas skyddshus
I Finland har vi fyra mycket olika årstider.
FPA:s kostnadsersättningfinska _ svenska _ engelska
Ring journumret 045 639 6274 om du behöver en plats på skyddshemmet.
linkkiMellersta Finlands tolkcentral:
Därefter ger TE-byrån ett utlåtande i ärendet till den instans som betalar förmånen, det vill säga till arbetslöshetskassan eller FPA.
Om du vill ha mera kunskap och färdigheter innan du söker till en yrkesinriktad utbildning, kan du ansöka till VALMA-utbildningen.
Också positiva saker, t.ex. att man får barn, kan ändra livet så mycket att man behöver stöd i den nya situationen.
Du kan få stöd för skolresor (koulumatkatuki) om du bor i Finland och studerar i gymnasiet eller vid en yrkesläroanstalt.
Fråga mer vid den läroanstalt där du vill studera.
Patientombudsmannens tjänster är kostnadsfria.
Om du är kund hos en mottagningscentral kan du ansöka om stöd för frivilligt återvändande vid din egen mottagningscentral.
Under samtalet får den som ringer hjälp med att kartlägga sin situation, råd och vid behov vägledning till något ställe där man kan få hjälp.
Rättighet
Som EU-medborgare behöver du inget arbetstillstånd i Finland.
Nybörjarnivån
Kontorets öppettider
Vad kan jag studera i yrkesinriktad arbetskraftsutbildning?
Privat dagvård och hemvårdsstöd
Observera att handlingarna ska vara på finska, svenska eller engelska.
Läs mer: Handikappade personer.
I Finland kan alla gifta sig som
I nödsituationer ringer du det allmänna nödnumret 112.
Du kan fråga vid närmaste FPA-byrå hur du kan få hjälpmedel.
Böcker och annat material finns på flera olika språk.
Om äktenskapet slutar i skilsmässa delas makarnas sammanlagda egendom jämnt mellan makarna.
Fyll i blanketten i Enter Finland-tjänsten.
Brott kan anmälas per telefon eller fax, på polisens webbplats eller genom personligt besök till polisstationen.
Service för missbrukarefinska _ svenska
Arbetsgivaren ska ge den anställda en skriftlig redogörelse för de centrala villkoren i arbetet vid tillsvidare gällande anställningar samt anställningar som varar över en månad.
Du kan resa till Finland om du har ett giltigt ID-kort eller pass.
hittar du en lista över webbsidor där du kan ansöka om bostad.
Uthyrning i andra hand
Läs mer på InfoFinlands sida Universitet.
registrerat uppehållstillstånd;
Läs mer: Trafik.
Rabatter för pensionärer
praktik projekt
Du ska ha med dig kortet på varje besök till rådgivningen.
Socialhandledare 016-322 3124, 040-729 8766
byta en säkring
Fackförbundets representant på arbetsplatsen
Till en del kurser kan du anmäla dig på Internet.
Du kan lära dig ett nytt yrke eller en ny examensdel.
Om en närstående dör oväntat och du behöver stöd kan du kontakta social- och krisjouren i Esbo, telefon (09) 816 42439.
För att barnet ska kunna få uppehållstillstånd måste hans/hennes uppehälle i Finland vara tryggat, till exempel genom förälderns löneinkomster.
Om du redan har finländsk personbeteckning och ett skattekort, hittar du skattenumret på ditt skattekort.
Tfn (09) 505 6379
Företagshälsovårdens tjänster
Den omfattar 12 kvarter med hundratals trähus och gårdsbyggnader.
tillräckliga kunskaper, färdigheter och resurser för den företagsverksamhet som du planerar
Att färdas på isen
Stöd vid skilsmässafinska
Vård av barnet
Teater och filmer
I det här fallet är tolkningen avgiftsfri. Tolkning ska alltid begäras i förväg.
Likväl utreds alla ansökningar som EU-medborgare skickar in.
Läs mer på InfoFinlands sida Diskriminering och rasism.
Du ska då bifoga till ansökan ett löneintyg för löner som du har fått.
Användningen av dem kan vara begränsad, men oftast är de öppna för alla.
Privata hälsovårdstjänster är dock avsevärt dyrare för kunden än offentliga.
Arbetsförmedlingstjänster
Stödboende för personer med psykisk ohälsa och missbruksproblemfinska
Ansökan till förskoleundervisningfinska _ svenska _ engelska
ränteavdrag på bostadslån
på ett daghem (päiväkoti)
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
Till exempel får syskon inte ha samma namn som första namn.
CV:t kan även vara en video, en portfölj eller en webbsida.
Enligt lagen i Finland måste arbetstagarna behandlas väl och de ska betalas lön.
Fundera på hur ditt kunnande motsvarar arbetsgivarens önskemål och krav.
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Underhållsbidrag för barn
Bostadssituationen varierar mycket mellan olika orter.
Öppningsoperationen gör förlossningen och undersökningarna under graviditeten lättare.
Du kan läsa mer om registreringen av modern på InfoFinlands sida Registrering som invånare.
Tolktjänster
En meritförteckning, eller ett CV, är en kortfattad och tydlig sammanfattning av ditt kunnande, din arbetserfarenhet och din utbildning.
Vaccinationer är en central del av förebyggandet av smittsamma sjukdomar hos barn. Barnrådgivningen ger barnet de vanliga vaccinationerna.
Sökandens livssituation och behov av understöd är ofta mycket olika.
Du får mer information om tolktjänsterna i din kommun på rådgivningen.
Gör en skriftlig anmälan till din arbetsgivare senast två månader innan du blir moderskapsledig.
Sexuellt våld
Invånarna i Esbo kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
äkta par och registrerade par sambor
Du får arbetslöshetsförmån under utbildningstiden.
linkkiEuropaskolan i Helsingfors:
Giltigt ID-kort eller pass
Läs mer på InfoFinlands sida Uppehållstillstånd för make eller maka.
Rasism (rasismi) innebär att man betraktar någon människogrupp eller en person som hör till gruppen som sämre än andra till exempel på grund av etniskt ursprung, hudfärg, nationalitet, kultur, modersmål eller religion.
Barnen äter tre måltider under dagen: frukost, lunch och mellanmål.
Om barnet inte är tryggt i sitt hem eller om situationen med barnet är mycket svårt, kan det fattas ett beslut om vård utom hemmet eller omhändertagande.
Om du inte har en hemkommun i Finland ska du be FPA utreda din rätt till den offentliga hälso- och sjukvården.
Yrkesubildning
Enkäterna är oftast på engelska, ibland även på andra språk.
Esbo huvudpolisstation
Mer information finns på Karleby kyrkliga samfällighets webbplats.
Arbetsgivaren kan t.ex. betala avgifter för en kurs i finska för din räkning.
Vård av barn Invånarparker och klubbar
Det är bra att inleda medicineringen så tidigt som möjligt.
Läroanstalten meddelar dig att du har antagits för studier med ett brev.
Hörselförbundet och Finlands Dövas Förbund är organisationer som arbetar för att förbättra hörselskadade personers ställning i samhället.
Du får studera i Finland högst 360 dagar när du gör en underrättelse om rörlighet.
Du kan också söka bostad via föreningen Suomen Opiskelija-asunto (Suomen Opiskelija-asunto) (SOA).
Följ väderleksrapporterna och använd alltid en flytväst i rätt storlek.
Du behöver intyget om du ansöker om moderskapsledighet av din arbetsgivare.
Användaren kan förhindra användningen av cookies i sina webbläsarinställningar.
När du har sökt asyl har du rätt att vistas i Finland medan din ansökan behandlas.
Föräldern kan då ha antingen ensam eller gemensam vårdnad om barnet.
Om dina inkomster blir mindre eller större under året, ska du beställa ett nytt skattekort.
Kontrollera regelbundet att brandvarnaren fungerar.
Om du flyttar utomlands för över ett år, betraktas flyttningen som permanent flyttning.
Eldstadsvägen 7 B, vån.
Hur du ringer nödnumretfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ arabiska _ kurdiska _ albanska _ tyska
Ansökan ska göras innan du har vistats utomlands över två år.
bedömningen av hur bra du kan klara av studierna.
Så här ansöker du om Schengenvisum
Det kallas för lättföretagande.
Möblerade hyresbostäder och lägenhetshotell
yrkesutbildning
via tjänsten Mina e-tjänster eller per telefon.
Arbets- och näringsbyrån anvisar invandrare till kurser i finska språket som ingår i integrationsprocessen.
Socialtjänsterfinska _ svenska _ engelska
Detta innebär att du håller en paus i lyftandet av pensionen.
Mer information om familjeåterförening finns på InfoFinlands sida Till familjemedlem i Finland.
I den inledande kartläggningen får du information om utbildning i finska eller svenska, arbetssökning, utbildning och tjänster i Vanda.
linkkiFöreningen för mental hälsa i Finland:
Ungefär fem procent av finländarna har svenska som modersmål.
Läs mer om finska medborgarnas rättigheter och skyldigheter på InfoFinlands sida Finskt medborgarskap.
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem (turvakoti).
Vandainfon finns i Dickursby, Korso och Myrbacka.
Anmälningstiden är i början av året, vanligen i januari.
Grundläggande utbildning
ABC för restaurangbranschen:
I Finland tillhandahåller kommunerna kommunal småbarnspedagogik bland annat i daghem.
När du söker sjukdagpenning ska du bifoga till ansökan:
Hemvårdsstödet består av en vårdpenning och ett vårdtillägg som är beroende av familjens inkomster samt ett eventuellt kommuntillägg.
Människorna samlas på picknick.
Fastställande av faderskap (Isyyden tunnustaminen)
linkkiInstitutet för hälsa och välfärd:
Du kan inte identifiera dig med ett körkort.
Också universitetet flyttades år 1828 från Åbo till Helsingfors.
Kurser – Lista kurserna i finska och andra kurser som du avlagt under en egen rubrik.
I Helsingfors finns det också privata skolor med undervisning på t.ex. engelska, tyska, franska eller ryska.
Från EES-länderna får du ta med dig den mängd läkemedel för eget bruk som motsvarar ett års förbrukning.
Även andra anhöriga till en person som har ett uppehållstillstånd på grund av internationellt skydd kan beviljas uppehållstillstånd.
Förtroendemannen väljs av de anställda.
en hyresbostad
Samtal på finska
Pensionsbeloppet beror på hur länge personen har bott eller arbetat i Finland.
Dit kallas brottsoffret, den brottsmisstänkta och vittnen.
Vissa preparat kan tas inom 120 timmar efter samlaget.
Du kan beviljas asyl i Finland om myndigheterna anser att du blir förföljd i ditt hemland på grund av
utan tvingande skäl göra upp öppen eld på annans mark
Ansökan till vissa universitetsstudier sker genom en separat ansökan.
Dessutom krävs det att du har haft din hemkommun i Finland i minst två år i rad.
Ingen får dömas till döden eller torteras.
En invandrarförening kan hjälpa dig att bevara och utveckla din kultur.
Familjerådgivningfinska _ svenska
Polska
Rättigheter
Umgängesrätten kan till exempel innebära att barnet bor hos den ena föräldern och träffar den andra föräldern vartannat veckoslut och dessutom vissa tider under loven.
Olika konstarter är musik, bildkonst, dans, teater, cirkuskonst, ordkonst, handarbete och arkitektur.
Om du har betalat för mycket i skatt, får du skatteåterbäring (veronpalautus).
Innan du skriver din jobbansökan, läs jobbannonsen noga och fundera på vilka färdigheter och vilket kunnande arbetsgivaren är ute efter.
Den har öppet dygnet runt.
Barn under 15 år behöver ett läkarrecept.
Bybibliotek linkkiBybiblioteken:
Kränkande eller osakligt innehåll
Med hjälp av gränssnittet kan du visa InfoFinlands innehåll på andra webbplatser eller skapa olika applikationer.
Traumatiska upplevelser
Information om tjänsterna finns på sidan Som invandrare i Vanda.
Fredrikinkatu 48
Helsingfors enhet
Hedersrelaterat våld kan vara till exempel
En del områden är väldigt populära. I sådana områden hyrs bostäderna ut mycket snabbt.
Tjänsterna vid A-kliniken i den egna kommunen är kostnadsfria för klienter som bor stadigvarande i Finland.
Regionala ungdomstjänsterfinska
I Helsingfors finns många privata läkarstationer som även tar hand om barn.
du ber en släktning eller vän gå i borgen för ditt lån.
Läs mer om vem som omfattas av den finländska sjukförsäkringen på InfoFinlands sida Den sociala tryggheten i Finland.
Malms sjukhus
Lapplands yrkeshögskolafinska _ engelska
Äldre människors hälsa.
Yrkeshögskolan kan ordna avgiftsfri utbildning för invandrare med målet att ge den studerande tillräckliga språkkunskaper och andra färdigheter som behövs för att studera vid yrkeshögskolan.
På InfoFinlands sida I Finland utan uppehållstillstånd finns det mer information för papperslösa.
Du kan få stöd om du på grund av ditt handikapp eller din sjukdom behöver kontinuerligt hjälp.
Tjänster för handikappadefinska
Privata hyresbostäder
Om du misstänker att ett barn har förgiftats kan du fråga råd vid Giftinformationscentralen (Myrkytystietokeskus).
Företagarens skyldigheter
För akutpreventivmedel behövs vanligen inget recept.
Problem i skolan eller med studierna
På gymnasiet behövs goda språkkunskaper.
Broschyren Att söka pension från utlandetfinska _ svenska _ engelska _ ryska _ estniska
pedagogiska områden
År 1946 inkorporerades nya områden till Helsingfors och staden yta mångfaldigades nästan åtta gånger.
Om du insjuknar plötsligt eller om du råkar ut för en olycka, får du akut sjukvård även om din hemkommun inte är Vanda.
Stämpeln ska begäras vid utrikesministeriet i det ifrågavarande landet och dessutom vid Finlands beskickning i landet.
Du kan ringa brottsofferjouren om du eller en närstående har blivit utsatt för ett brott eller om du har bevittnat ett brott.
Telefonrådgivning: (09) 816 45285
arbetsgivarens och arbetstagarens hemort eller driftställe
Karleby handelsflotta var under perioder Finlands största.
Ekonomi- och skuldrådgivning ordnas av kommuner.
Ett försäkringsintyg eller en kopia av det europeiska sjukvårdskortet
MoniNet är ett mångkulturellt center i Rovaniemi, Lappland.
Rådgivningsbyrån för familjeplanering ger stöd i frågor om familjeplanering och graviditetsprevention.
Stöd till företagare
Du får information om hur du köper läkemedel på InfoFinlands sida Läkemedel.
Arbetsgivaren måste följa kollektivavtalet.
Information om hälsorådgivningfinska _ svenska _ engelska
Rådgivningen betjänar telefonledes på numret 045-237 7104 (måndagar kl. 14–16).
Naturens husfinska _ svenska _ engelska
linkkiVanda stad:
På samma adress ser du också hur behandlingen av din ansökan framskrider.
Om du till exempel orsakar en vattenskada måste du själv betala hela renoveringskostnaden.
I studiemiljön finns sju avsnitt som handlar om invandrarens liv i Finland.
Vilka reklammedel ska du använda för att främja försäljningen?
Rehabiliteringsstöd är invaliditetspension på viss tid.
Läs mer: Fortsatt uppehållstillstånd.
I Karleby är den kemiska industrin och industri i anslutning till denna särskilt viktig.
Erkännande (BY) – Du måste nämna källan InfoFinland.fi.
I nödsituationer ringer du nödnumret 112.
När arbetsavtalet gäller tillsvidare har arbetstagaren en fast eller permanent anställning.
För fristående yrkesexamen finns ingen bestämd ansökningstid.
Vad händer i småbarnspedagogiken?
Ibland kan norrsken ses också i södra Finland.
registrerad partner
Enligt Finlands lag ska hinder mot äktenskap prövas om du är finsk medborgare eller permanent bosatt i Finland och uppgifterna om dig finns i befolkningsregistret.
Man kan dock använda bilen tillfälligt innan bilskatten är betald.
I Finland finns många medborgarinstitut (kansalaisopisto) och arbetarinstitut (työväenopisto).
Skolhälsovårdfinska _ svenska
I Helsingfors finns såväl universitet som yrkeshögskolor.
Bouppteckningen ordnas av den person som bäst känner till den avlidnes egendom och skulder.
direkt via lönesystemet om det har en inbyggd teknisk förbindelse till Inkomstregistret eller
Läs mer på InfoFinlands sida Till familjemedlem i Finland.
När perioden har gått kan man ansöka om förlängning för bidraget.
Den förberedande undervisningen varar vanligtvis ett år.
På stadens webbplats hittar du kontaktuppgifterna till skolorna och mer information om anmälan.
I vissa enskilda fall kan man avvika från försörjningsförutsättningen om det finns exceptionellt vägande skäl eller om barnets bästa kräver detta.
Hjälp med att få slut på våld
Läs mer om barndagvård, förskoleundervisning och grundläggande utbildning på InfoFinlands sida Utbildning för barn.
Man måste delta i rättegången.
Du måste ansöka om familjeförmåner separat från FPA.
Motion och friluftsliv i Helsingforsfinska _ svenska _ engelska
Sambor kan även upprätta ett skriftligt avtal om hur egendomen ska fördelas om paret går isär.
Om du är medborgare i ett EU-land, Liechtenstein eller Schweiz och vill resa till Finland för en kort period, till exempel på semester, på affärsresa eller för att besöka släktingar, behöver du inget visum.
Läs mer: Tandvård.
I Finland är det vanligt med familjer med en förälder.
02700 Grankulla
Tolkningfinska _ svenska _ engelska
Du kan utnyttja de offentliga hälsovårdstjänsterna i Finland om du har hemkommun (kotikunta) i Finland.
Du kan också leta upp en privat familjedagvårdare som vårdar barnen hemma hos sig, eller anställa en skötare i ditt eget hem.
Du kan också hämta ansökningsblanketten på daghemmet eller vid informationen i stadshuset.
Arbets- och näringsbyråerna i Nylandfinska _ svenska
reparera en enfas skarvsladd (spänning 230 V)
Information om det europeiska sjukvårdskortetfinska _ svenska _ engelska
gymnasiet
Begravningstillstånd
EU-medborgarnas rättigheter som rätten att fritt röra sig och arbeta inom EU:s område och rätten att rösta och ställa upp som kandidat i EU-val
Även kommunerna äger hyresbostäder. De är ofta förmånligare än andra hyresbostäder.
Telefonnumret till den gemensamma telefontjänsten för hälsostationerna i Vanda är 09 839 50 000.
Grundskoleelever får stöd i sitt skolarbete.
Stöd för frivilligt återvändandefinska _ svenska _ engelska _ persiska _ arabiska
Broschyren Makens efternamn och barnets efternamnfinska _ svenska _ engelska
Adjektiven böjs efter dessa genus.
Du kan be om att få tid hos en kvinnlig läkare om du vill.
Besök läkaren före slutet av den fjärde graviditetsmånaden.
I Finland råder religionsfrihet.
Om dina studier i Finland till exempel varar mindre än två år, ska försäkringen täcka sjukvårdskostnader upp till minst 100 000 euro.
Studietiden beror på utbildningsprogrammet och din egen studietakt.
Sysselsättningsutsikter för olika yrken i Finlandfinska _ svenska _ engelska
Det är bra att beakta att parförhållandets form påverkar makarnas rättigheter och skyldigheter, frågor som rör egendom och arv, vårdnad om och underhåll av barn samt adoption.
Den lön som betalas till arbetstagaren är nettolönen (nettopalkka).
Finlands Röda Kors hjälper med att ordna resan till Finland för kvotflyktingens familjemedlemmar när dessa fått uppehållstillstånd.
Du kan diskutera preventivmetoder med skolans hälsovårdare och i vissa kommuner kan skolans hälsovårdare ge dig ett startpaket.
Fråga mer hos FPA.
När du ansöker om en förmån, utreder FPA om du har rätt till FPA:s förmåner.
I vuxenutbildningen avlägger du yrkesexamen som fristående examen.
hittar en arbetsplats eller studieplats,
Du kan också söka till ett separat magisterprogram.
linkkiHälsovårdscentralen:
Du får anvisningar om hur detta påverkar ditt utkomststöd för arbetslösa.
I norra Finland kan temperaturen vara till och med -30 grader.
Mer information om att ansöka om skilsmässa hittar du på justitieministeriets webbplats.
Skolbyrån
För att arbeta måste du ha ett finländskt skattekort.
Du ska ansöka om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut.
Boka tiden via Migrationsverkets elektroniska tidsbokningssystem.
Läs mer om utlänningars rösträtt i Finland på InfoFinlands sida Val i Finland.
I Vanda finns även Finavia Avia College som ger utbildning för olika luftfartsyrken.
Integrationsutbildningen kan omfatta studier i finska, andra studier eller arbetsförsök.
Ansökan om ordningsnummerfinska _ svenska _ engelska
Till exempel FPA och migrationsverket (Maahanmuuttovirasto) beställer i vissa fall en tolk för kunden.
EU-medborgare ska också registrera sig på Migrationsverket.
linkkiEsbo biIdkonstskola:
Om du har problem med alkohol eller andra droger eller spelproblem kan du ta kontakt med A-klinikkaan.
Du kan samtidigt köpa fler andelar i din bostad om du har kommit överens med byggherren om detta.
Preventivrådgivningfinska _ svenska _ engelska
linkkiPyhäjoki kommun:
Reseplanerarefinska _ svenska _ engelska _ ryska
Serviceboendefinska _ svenska _ engelska
Det är möjligt att i enskilda fall avvika från försörjningsförutsättningen, om det finns exceptionellt vägande skäl eller om barnets bästa kräver detta.
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en krismottagning för invandrare.
Boendetiden kan vara från en dag till flera månader.
Information om Finland till turistersvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Då hyrsvärden väljer hyresgäst får han eller hon enligt lagen inte diskriminera någon exempelvis på grund av etniskt ursprung, religion eller nationalitet.
Besök Migrationsverkets tjänsteställe; du måste styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Alla invandrare har rätt att få grundläggande information om Finland.
Förberedande utbildning för invandrare
Blivande förskolebarn får mer information om detta per post, på dagvårdens webbplats och i lokaltidningen.
Tandvården vid hälsovårdscentralen är avgiftsfri för barn under 18 år.
Läs mer på InfoFinlands sida Våld och Hedersrelaterat våld.
Röda Korset söker försvunna anhöriga och förmedlar meddelanden på krisområden.
Det är inte obligatoriskt att ta studielån.
Därefter kan man fortsätta studierna och avlägga yrkesexamen eller specialyrkesexamen.
I Finland finns också slott som är öppna för allmänheten, till exempel Olofsborg, Åbo slott och Tavastehus slott.
Vanligtvis ansöker man om dagvårdsplats i den egna kommunen.
Deras färdighetsnivå är 1–2.
Naturen i Finland är mångsidig.
Gifta makar av samma kön har rätt att adoptera ett barn och rätt till adoption inom familjen.
Du kan även be om hjälp och råd vid kommunens skuldrådgivning eller socialverk eller en boenderådgivare vid kommunen eller hyreshusbolaget eller till exempel Garantistiftelsen.
Uppehållstillstånd på andra grunderfinska _ svenska _ engelska
Med den här blanketten kan du meddela följande information till myndigheterna:
linkkiEuropeiska unionen:
Svenska språket i Finland.
Var ligger närmaste magistrat, hälsostation eller bibliotek?
Distansgymnasiumfinska
När du flyttar i Finland från en bostad till en annan:
Information om tågtidtabellerna hittar du på VR:s webbplats och på järnvägsstationerna.
När hemvården är regelbunden påverkar dina egna och din makas eller makes inkomster hemvårdsavgiften.
Broschyren Information till asylsökandefinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Läs mer om att bevisa dina språkkunskaper på InfoFinlands sida Officiellt intyg över språkkunskaper.
I Helsingfors finns det flera daghem som drivs av staden och privata daghem.
Motion
Samtalen besvaras av krisarbetare och utbildade frivilliga stödpersoner.
I Finland värdesätts ärlighet.
Fyll i blanketten noggrant och underteckna den.
Då är barnet ca nio månader gammalt.
Om umgänget blir problematiskt
Färdighetsnivåerna i statsförvaltningens språkexaminafinska _ svenska
Rasism och rasistiska brott
Om föräldrarna är gifta kan de välja endera makens efternamn till barnet.
I krissituationer kan du ringa eller åka till jouren.
Ett samboförhållande registreras inte någonstans.
Film om munhälsovårdfinska _ engelska _ somaliska _ arabiska
Läs mer på InfoFinlands sida Rättigheter och skyldigheter för boende.
Tfn (09) 816 45285
till vård av hög kvalitet
Rådgivningen ges av en jurist.
Asylsökande
linkkiMellersta Österbottens social- och hälsovårdssamkommun Soite:
En rörelsenedsättning kan bero på en sjukdom, ett olycksfall eller genetiska orsaker.
Vård utom hemmet betyder att barnet bor någon annanstans än hos sina föräldrar.
Ryska och engelska: 050 325 7173
I ett höghus hittar du ordningsreglerna vanligtvis i trapphuset nära entrédörren.
Om du vistas i Finland utan uppehållstillstånd kan du emellertid bli tvungen att betala för vården.
Vad stadigvarande boende betyder definieras i lagen.
Sambo med en utländsk medborgare
Alla helgons dag firas i början av november.
linkkiKommunbostäder:
Fundera på vilka produktionsmedel eller vilken arbetskraft du behöver.
Mer information om den kommunala ungdomsverksamheten får du hos ungdomsväsendet i din hemkommun.
Ibland finns det i annonsen en utsatt tid då bostaden visas.
Studietillfällena är dock öppna för alla.
Vad är våld?
arbete
När du flyttar ditt stadigvarande boende till Helsingfors, ska du registrera dig som invånare i kommunen.
Ansökan ska lämnas in till FPA senast en månad innan moderskapspenningperiodens utgång och föräldrapenningperiodens början.
Karlebygatan 27, PB 581
Sambor kan ha sådan egendom om vars ägande de inte har en överenskommelse.
linkkiFinansministeriet:
Stadsfullmäktiges sammanträden på Internetfinska
Medborgarinstitutens musikgrupper är öppna för alla.
Bouppteckningshandlingen (perukirja) ska lämnas till skattebyrån senast en månad efter bouppteckningen.
Prövningen tar ungefär en vecka.
Om du söker till ett utbildningsprogram där undervisningsspråket är ett annat än finska eller svenska, beror ansökningssättet på utbildningen.
Boka en tid hos hälsostationens allmänläkare om du till exempel har problem med blödningar eller smärtor i underlivet.
eBiblioteket (eKirjasto) tillhandahåller elektroniska material, såsom böcker, tidskrifter och filmer.
På babyresa - För dig som har fött barnfinska _ svenska _ engelska
Om du har problem eller oklarheter med uppehållstillståndet, kan du ta kontakt med följande instanser för att be om råd:
Du kan bli klient om du flyttat till Finland på grund av familjeband, är flykting, offer för människohandel eller har rätt till en inledande kartläggning.
Vanligtvis är barnets föräldrar dess vårdnadshavare.
Information om skolresestödetfinska _ svenska _ engelska
När du funderar på vilken företagsform du ska välja, är det absolut tillrådligt att du kontaktar företagsrådgivningen.
–15 studeranden och vanligtvis finns det 8–10 undervisningsgrupper.
Fackets ABC-bokfinska _ engelska _ ryska _ estniska
Fråga mer vid din läroanstalt.
Yrkesexamen och specialyrkesexamen ger dig behörighet till ett visst yrke.
Den förberedande utbildningen tar ett läsår och ger beredskap för gymnasiestudier.
som har rösträtt i val till Europaparlamentet och
Information om fackförbundsverksamhetfinska _ svenska _ engelska
I naturhuset Villa Elfvik ordnas utflykter, evenemang och utställningar.
Tfn (09) 5056 357 eller (09) 5056 358
Ateneumfinska _ svenska _ engelska
Broschyren Information om den finska grundskolanengelska _ ryska _ franska _ somaliska _ arabiska
Religiösa seder eller ritualer hör inte hemma på den finländska arbetsplatsen.
Samtidigt får du en ansökningsblankett.
Som bevis duger till exempel ett utdrag ur boenderegistret eller ett hyreskontrakt med bådas namn.
hushållets bruttoinkomster (inkomster före skatt)
Det är bra att ni går till kliniken tillsammans.
Om det behövs kan du få servicerådgivning om användningen av nättjänsterna.
Söndagen är påskdagen och då minns man Jesu uppståndelse.
Ta reda på om du kan skjuta upp andra betalningar för att kunna betala hyran.
Livet kan vara svårt till exempel när man flyttar från ett land till ett annat, har problem på arbetsplatsen, förlorar sin arbetsplats, har problem i familjen, går igenom skilsmässa, förlorar en anhörig, blir sjuk eller när livet förändras på andra sätt.
Mer information hittar du på Helsingfors stads webbplats.
Via tjänsten Religionerna i Finland kan du söka information enligt religionssamfund och ort.
I Helsingfors har papperslösa invandrare rätt att få brådskande och nödvändig vård inom de offentliga hälsovårdstjänsterna.
Kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
Borgerliga vigslar förrättas på magistraten.
Du kan få fortbildning eller påbyggnadsutbildning i din egen bransch.
Tfn 045 639 6274 (24h)
Flyttanmälanfinska _ svenska _ engelska
Barnet får utföra lätt arbete några timmar om dagen om det inte skadar hennes hälsa eller skolgång.
linkkiRättsväsendet:
linkkiAnonyma alkoholister, AA:
Yrkesexamen kan även avläggas med läroavtal.
Företagshälsovård
Hur du ansöker om pension till utlandet beror på i vilket land du bor.
Behöver jag ett tillstånd för företaget?
Tjänster av detta slag är bland annat måltidstjänst och transporttjänst.
Du kan delta i yrkesinriktad arbetskraftsutbildning, om
Studerandena inom integrationsutbildningen kommer från tiotals olika länder och undervisningsspråket är finska. En kurs kan ha 8
I dagvården lär barnet känna den finländska kulturen, lär sig det finska språket och verkar i en social grupp.
Längst ner på varje undersida i InfoFinland hittar du en responslänk, via vilken du kan skicka respons som direkt berör innehållet på sidan.
Vård av barnet i hemmet
17 år
Också många arbetsplatser utbildar sina anställda till exempel i användningen av nya apparater eller program.
Om du flyttar ditt stadigvarande boende till Grankulla, ska du registrera dig som invånare i kommunen.
Läroplikten upphör om den inte redan har fullgjorts.
Vasavägen 7
Du måste ansöka om ett nytt uppehållstillstånd på grund av arbete innan ditt uppehållstillstånd för att söka arbete går ut.
Vid Vanda vuxenutbildningsinstitut (Vantaan Aikuisopisto) kan man till exempel skapa konst, handarbeten, laga mat eller dansa.
Om du har en sjukförsäkring i ett annat EU-land, EES-land eller i Schweiz har du rätt till nödvändig sjukvård i Finland.
Vid folkhögskolor kan du även avlägga yrkesexamen.
Rätten till FPA:s förmåner
Böle verksamhetsställe
Fråga bibliotekarienfinska _ svenska _ engelska
Enligt lag har du rätt att välja antingen finska eller svenska som integrationsspråk.
Vissa tv-program kan du titta på avgiftsfritt.
Avdragen beaktas då i din skatteprocent.
Bibliotek
En del arbetsgivare utbildar människor till arbeten hos dem.
Om studeranden har ett annat modersmål än finska eller svenska och saknar tillräckliga språkkunskaper för gymnasiestudierna, kan hen söka till förberedande gymnasieutbildning (LUVA).
Söka tjänster
Merparten av studierna är dock på finska eller på svenska.
linkkiMiljöförvaltningen:
Välkommen!
Utbildning för döva invandrarefinska _ svenska _ engelska
Du kan studera finska som arbetskraftsutbildning.
Den förberedande undervisningen före grundskolan är avsedd för alla de barn med invandrarbakgrund som inte har tillräckliga kunskaper för att klara sig i undervisningen inom den grundläggande utbildningen.
Du själv betalar förmedlingsarvodet endast om du har ingått ett skriftligt uppdragsavtal med bostadsförmedlaren om att söka en bostad åt dig.
På universitet kan man avlägga lägre högskoleexamen på cirka tre år och därefter högre högskoleexamen på cirka två år.
Läs mer: Läkemedel.
Uppehållstillstånd för arbetstagare
handikappade
Mer information om den allmänna språkexamen får du på Utbildningsstyrelsens webbplats.
Om du har fyllt 61 år kan du få partiell pension redan före din lägsta ålderspensionsålder.
Integrationscentret Kotoutumiskeskus Monika hjälper arbetslösa invandrarkvinnor att hitta jobb.
Lämna in ansökan till daghemmet eller stadshuset.
dagvård
Då måste du betala för operationen själv.
Övriga hyresbostäder
Fackförbundets medlemmar betalar förbundet en medlemsavgift som vanligen är cirka 1–2 procent av lönen.
Nödnumret (hätänumero) i Finland är 112.
Målsättningen med verksamheten är att främja barnets utveckling och lärande.
Om du har uppehållstillstånd och hemkommun i Finland, har du rätt till kommunens tjänster för handikappade.
Vi svarar på responsen på följande språk: finska, svenska och engelska.
Meddela din arbetsgivare om familjeledigheten senast två månader innan den börjar.
Diagram över erkännande av examen(pdf, 410,87 kt)finska _ svenska _ engelska
Arbets- och näringsbyrån genomför utbildningar även tillsammans med arbetsgivare.
Om du är berättigad till integrationsstöd ska du kontakta TE-byrån innan du ansöker.
På MoniNets webbplats finns länkar till olika webbsidor där du kan studera finska på egen hand.
Ibland inleds förlossningen normalt men akut kejsarsnitt blir nödvändigt på grund av barnets tillstånd.
Fråga bibliotekarien-tjänsten
Offentlig rättshjälp söks vid statens rättshjälpsbyråer.
Efter betänketiden fullföljer man sin ansökan med en ny ansökan.
att vid behov få hjälp av patientombudsmannen (potilasasiamies).
Då har du inte rätt till FPA:s förmåner.
Du kan betala för taxin med kontanter eller med bank- eller kreditkort.
Läs mer om frivilligarbete på InfoFinlands sida Frivilligarbete.
Om du inte behöver brådskande tandvård, ring efter kl. 10.00.
Ranunkelvägen 22
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Möten måste avtalas på förhand.
Mentalvårdsenheterna har verksamhet på två adresser:
antalet vuxna och barn i hushållets storlek
Brådskande fall sköts så fort som möjligt.
Om någon bryter in sig i ditt hem, ring nödnumret 112.
modern har en hemkommun i Finland och
Barnbidragsbeloppet är en aning högre för varje följande barn.
Om du nyligen har flyttat till Finland, måste du registrera dig som invånare.
I Finland är det vanligt att köpa använda saker och lätt att hitta använda saker i gott skick.
Om du har en långvarig sjukdom ska du ta med dina gamla recept till läkarmottagningen så kan läkaren beakta dessa när han eller hon skriver ut ett recept.
Den tryckta guiden finns i företagsservicecentralerna i kommunerna på området.
föräldradagpenning
Läs mer på InfoFinlands sida Beskattning.
Västra Nylands rättshjälpsbyrå
Kommunalval
linkkiMannerheims Barnskyddsförbund rf:
Du kan även ta kontakt på en annan persons eller på någon grupps vägnar.
Information om jämställdhet i arbetslivetfinska _ svenska _ engelska _ ryska _ samiska
Från Rovaniemi flygplats finns flera flyg till Helsingfors, andra städer i landet och utrikes resmål.
Tjänsterna kan variera något i olika delar av landet.
Om ett invandrarbarn går i en skola där undervisningsspråket är finska studerar barnet också svenska som främmande språk tillsammans med de finskspråkiga eleverna.
i ett privat daghem eller i ett gruppfamiljedaghem
linkkiArbets- och näringsbyrån:
ange exakt adress och kommun
Om du har ingått äktenskap med en finländsk medborgare som är bosatt i Finland kan du få uppehållstillstånd i Finland på grund av familjeband.
Yle är en offentlig tjänst och dess verksamhet bekostas med skattepengar.
Ange i slutet av videoklippet namnen på samtliga personer som medverkat i skapandet av videoklippet.
Problem med uppehållstillstånd
Också ett barn till utländska föräldrar som föds i Finland kan få finskt medborgarskap, om hen inte får medborgarskap i något annat land av sina föräldrar.
Man kan få ett flerårigt fängelsestraff för det.
Arbetspensionsutdraget visar hur stor pension du tjänat in i Finland.
Om en annan vårdnadshavare än barnets mor eller far ansöker om uppehållstillstånd måste vårdnaden bevisas till exempel genom uppvisande av ett domstolsbeslut.
Om du avser ansöka om startpenning ska du kontakta arbets- och näringsbyrån i ett så tidigt skede som möjligt.
Du hittar mer information om världsarven på Museiverkets webbplats.
Det är bra att reservera tid för detta eftersom förfaringssätten varierar i olika länder.
Om du ansöker om en dagvårdsplats i stadens daghem, ska du skicka in din ansökan minst fyra månader före dagvårdsstart.
Det är bra att skriva upp felen i bostaden tillsammans med hyresvärden när hyresförhållandet inleds.
Beskickningarna hjälper sitt lands medborgare som hamnat i nödläge i Finland.
Det är vanligt att par lever i ett samboförhållande före äktenskapet.
Vanda stads tjänster för invandrare omfattar
Du kan anmäla ditt barn till skolan i närskolan.
Mer information och anmälan finns på NewCo Helsinkis webbplats.
Tåg
Nöteborgsfreden 1323 avslutade kriget mellan Sverige och Novgorod om herraväldet i området.
Kontaktuppgifter till privata läkarstationer hittar du till exempel på internet.
du behöver startpengen för ditt uppehälle
Du kan få rehabiliteringspenning på samma villkor också när din hemkommun ordnar din rehabilitering.
Om du har en gammal tv, behöver du också en digitalbox för att titta på tv-program.
med en allmän språkexamen (yleinen kielitutkinto)
Fundera på hur du ska lyfta fram ditt kunnande och din lämplighet för uppgiften.
När du öppnar ett bankkonto lönar det sig att även skaffa webbankkoder.
I de flesta utbildningsprogrammen är undervisningsspråket ändå finska eller svenska.
Tolkning vid förlossningen
När äktenskapet slutar kan ni gemensamt komma överens om hur ni delar egendomen.
Social- och krisjourenfinska _ svenska _ engelska
Om hen inte kan hjälpa dig, ska du kontakta arbetsplatsens arbetarskyddsfullmäktige eller förtroendeman.
Lapplands yrkeshögskola
I Helsingfors kan du avlägga högskolestudier i många branscher.
Om man deltar i möten kan man påverka, föreslå ändringar och utveckla sitt eget arbete.
Chatten betjänar på finska, engelska, ryska och arabiska.
Vissa kommuner erbjuder unga kostnadsfria preventivmedel.
är 22 år gammal, har medborgarskap också i en annan stat och saknar tillräcklig anknytning till Finland
Finland har varit bebott sedan istiden, från cirka år 8800 före tideräkningen.
Om du är studerande kan du ansöka om en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS (Helsingin seudun Opiskelija-asuntosäätiö HOAS).
Motion för handikappade barn och ungafinska _ svenska _ engelska
Arbetsplatser i kommunernafinska _ svenska _ engelska
Läs mer på InfoFinlands sida Flytta från Finland.
Riksdagsval förrättas vart fjärde år.
Det är avgiftsfritt att delta i grupperna.
Grundläggande information om fortbildningfinska _ svenska
Också din arbetsgivare kan göra anmälan.
Priser på hyresbostäder med statliga stödengelska
För den som flyttar till Finland är det viktigt att känna till de grundläggande reglerna som gäller i arbetslivet och det finländska samhället.
Man kan till exempel prata om barnens situation i medlingen.
Medborgare i alla länder kan gifta sig i Finland.
Äkta makar är sinsemellan likvärdiga.
På hälsostationerna finns vanligtvis läkarens, sjukskötarens och hälsovårdarens mottagningar.
Registreringen kan göras till exempel på besiktningsstationer, vid försäkringsbolag och hos bilhandlare.
Kom ihåg att ansöka om särskild moderskapspenning hos FPA inom fyra månader från den dag du slutar arbeta.
Företagsfinland (Yritys-Suomi) (webbplats och telefontjänst)
Vanligen vårdar någondera av föräldrarna barnet i hemmet åtminstone under föräldraledigheten, det vill säga tills barnet är ca 9 månader gammalt.
Handläggningstider för tillståndsansökningarfinska _ svenska _ engelska
Barnet kan ha finskt medborgarskap och medborgarskap i något annat land.
Stadens hyresbostäder är vanligtvis förmånligare än de bostäder som hyrs ut av företag och privatpersoner.
profilområden: forskning i arktiska och nordliga frågor och forskning inom turism.
Läs mer om bostadsbidrag för sambor på InfoFinlands sida Bostadsbidrag.
Finland som en del av Kejsardömet Ryssland 1809–1917
Invalidpension betalas till 16–64-åringar.
Information om integration på svenskafinska _ svenska
Vid Lapplands yrkesinstitut kan du studera och skaffa dig yrkesinriktad grundutbildning och vuxenutbildning i alla studieområden förutom inom idrottsområdet och turism-, kosthålls- och ekonomibranschen.
På grund av ditt handikapp kan du även få rabatt på kollektivtrafikens biljettpriser.
Du kan fakturera vi en faktureringstjänst utan att starta ett eget företag.
Detta belopp påverkar inte ditt bostadsbidrag.
Efter lågkonjunkturen uppstod det mycket högteknologisk industri och högteknologiska arbetsplatser i Finland.
att göra en anmärkning till den vårdande enheten om patienten är missnöjd
På några orter finns det dessutom ledd motion som är avsedd endast för invandrare, exempelvis egna grupper för kvinnor eller för personer som vill bekanta sig med nya idrottsgrenar.
Yrkesexamen (ammattitutkinto)
Du kan bli kund vid Kompetenscentret via TE-byrån eller social -eller hälsovårdsverket.
Du kan söka till en yrkeshögskola för att avlägga en yrkeshögskoleexamen, då du har avlagt t.ex. någon av följande utbildningar:
Vanda stads hyresbostäder ägs och hyrs ut av VAV Asunnot Oy.
Detta kallas förvärvsinkomstavdrag (ansiotulovähennys).
Du kan gå till akutmottagningen vid akuta sjukfall där du inte kan vänta till följande dag på vård. Sådana fall är till exempel blödande sår, bröstsmärtor, brännskador med mera.
Då avfallet sorteras rätt kan man använda materialet för att tillverka nya produkter.
I stadsfullmäktige sitter 67 ledamöter som representerar olika politiska grupper.
Du kan även fråga om råd vid Helsinki-info.
På InfoFinlands sida Problem i äktenskap och parförhållande hittar du information om var du kan söka hjälp för problem i förhållandet.
Du kan också fråga om din egen situation vid FPA:s kontor eller telefontjänst.
Utvecklingsstörningen upptäcks ofta i barndomen eller ungdomen.
Om jämlikhet i arbetslivet föreskrivs i lagen om likabehandling och i arbetsavtalslagen.
Det är lätt att på ett pålitligt sätt hitta väsentlig information om integration av invandrare och om att bo i Finland på ett ställe, www.infofinland.fi.
Innan du besöker magistraten kan du fylla i Registreringsanmälan för utlänningar som finns på adressen maistraatti.fi.
Kontaktuppgifterna till vuxengymnasierna finns på Helsingfors stads webbplats.
Centrumbiblioteket Oodi, adress: Tölöviksgatan 4
15 år
Karlebys historiafinska _ svenska _ engelska
Riksomfattande kristelefonfinska _ svenska _ engelska
Läs mer: Hälsovårdstjänster i Finland
Ett kompetensbaserat CV lyfter fram ditt kunnande, dina färdigheter och dina erfarenheter.
Att hyra ut en del av bostaden till en annan person, om detta inte medför olägenhet för hyresvärden.
Då kan du söka direkt till läroverket i den separata ansökningsprocessen som är avsedd för dem som redan avlagt examen.
Hyresvärdar och banker kontrollerar ofta kredituppgifterna i kreditupplysningsregistret.
Läs mer om grunderna för uppehållstillstånd i InfoFinlands avsnitt Icke EU-medborgare.
Information om motionstjänsternafinska _ svenska _ engelska
Att bo i hyreslägenheten enligt vad som anges i hyresavtalet.
I avtalet ska den regelbundna arbetstiden nedtecknas.
linkkiFlyktinghjälp:
Riksomfattande kristelefon: 010 195 202
Genom att själv följa med arbetspensionsutdragen kan du kontrollera att din intjänade pension räknats rätt.
Joensuu
utvecklingsstörda
Läs mer:Vård av barnet.
Vårdnadshavaren måste underteckna arbetsavtalet.
Olika instanser ordnar företagarkurser och informationsmöten som är mycket nyttiga för dig som ska grunda ett företag.
Rovala 5
Lediga tjänster vid Esbo stad hittar du på stadens webbplats.
Föreningar bedriver sin verksamhet vanligen ett år i taget.
Enligt dessa ska anställda behandlas lika när det gäller anställning, arbetsförhållanden, anställningsvillkor, utbildning för personalen och avancemang i karriären.
Ta kontakt med TE-byrån så tidigt som möjligt om du ämnar ansöka om startpeng.
Tfn (09) 8392 4005
Du kan ansöka om en plats i stadens barnklubbar med blanketten som finns på stadens webbplats.
Fpa betalar barnförhöjningen tills barnet fyller 16 år.
Information för viseringsfria personer
Dagvård
barnet har någon annan privat skötare.
I vissa fall ersätter Kela en liten del av kostnaderna för privat sjukvård.
Skyddshemmen har jourmottagning dygnet runt.
I vissa städer får du använda tjänsterna vid mödrarådgivningen även om du vistas i Finland utan uppehållstillstånd.
Barnskyddslagenfinska _ svenska _ engelska
Hur står det till?
Du får bo i en bostadsrättsbostad om du först betalar bostadsrättsavgiften (asumisoikeusmaksu).
Tfn (09) 50 561
Studiernas omfattning är 60 eller 90 studiepoäng.
Ansökningstiden är i januari, men ansökan kan även lämnas in övriga tider, om familjen till exempel flyttar till Vanda mitt under året.
Det är möjligt att få en plats snabbare om den behövs för att du exempelvis erhållit arbete eller studieplats.
Om du inte kan betala din hyra
Om föräldrarna inte är överens, kan modern fatta beslut om religionstillhörigheten för ett barn som inte har fyllt ett år.
Besök läkaren vid rådgivningsbyrån före slutet av den fjärde graviditetsmånaden.
Arbetsgivaren ska ha en välgrundad orsak för att säga upp en anställd.
Finska medborgare har utöver det ovan nämnda också några ytterligare rättigheter och skyldigheter som utlänningar bosatta i Finland inte har.
Partiell sjukdagpenning ska sökas inom två månader efter att du börjar arbeta på deltid.
Långvarig sjukdom och vård av ett handikappat barn
Infobankens redaktion utser tävlingens vinnare i samråd med Infobankens användarråd.
Finland och Sovjetunionen ingick 1948 ett avtal om vänskap, samarbete och bistånd, enligt vilket staterna lovade att försvara varandra mot yttre hot.
I livshotande situationer ska du ringa nödnumret 112.
Böle verksamhetsställe
Läs mer:
Läs mera på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
Uppstartsföretagare
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
På InfoFinlands sida Arbetstagare eller företagare finns mer information för arbetstagare som flyttar till Finland.
bostadsbidrag för pensionstagare
Du kan ringa detta nummer om du behöver rådgivning i behandlingen av en sjukdom eller vill boka eller avboka en läkartid.
Barn får till exempel inte slås eller luggas.
Familjemedlemmarnas underhållsskyldighet sträcker sig inte till släktingar, till exempel vuxna syskon eller mor- eller farföräldrar.
På FPA:s webbplats finns en räknare som du kan använda för att beräkna om du uppfyller arbetsvillkoret för företagare.
Intyget över hindersprövningen ska finnas med vid vigselförrättningen.
Hälsotillståndet hos barn under skolåldern följs i barnrådgivningen (lastenneuvola).
Alla stater godkänner dock inte flerfaldigt medborgarskap.
Karleby är en teaterstad med långa anor, som erbjuder scenkonst på hög nivå framförd av både proffs och amatörer.
Information om dessa hittar du på webbplatserna för Informationscentralen för teater i Finland på finska, svenska och på engelska.
Den öppna linjen betjänar på finska, svenska och engelska.
Särskilt stöd erbjuds barn med handikapp inom småbarnspedagogiken och skolan.
Det samhällsvetenskapliga, företagsekonomiska och administrativa området
Onödiga samtal kan orsaka att hjälpen kommer för sent i verkliga nödsituationer.
Du kan också fråga om möjligheterna till rehabilitering, studier, arbete och hobbyer.
Du får vård på samma villkor och till samma kostnad som finländarna.
Om inkomsterna är mycket låga bortfaller bassjälvrisken.
Kom även ihåg att en underskrift är ett bindande avtal. Läs noga igenom alla dokument innan du undertecknar något.
Arbets- och näringsbyrån (TE-toimisto) kan hjälpa dig att hitta ett jobb.
Arbetsgivaren är också skyldig att göra de anställda förtrogna med arbetsplatsens säkerhetsanvisningar och lära dem korrekta arbetssätt.
Om du har hemkommun i Finland kan du ansöka om flexibel vårdpenning (joustava hoitoraha) för vård av barn under tre år och partiell vårdpenning (osittainen hoitoraha) för vård av skolbarn i årskurserna 1 eller 2 hos FPA.
Migrationsverket utreder din identitet och resväg till Finland och bedömer om du kan beviljas asyl i Finland.
linkkiFimea:
Till exempel motsvarar statsförvaltningens språkexamen som gäller goda språkkunskaper ett mognadsprov (kypsyysnäyte) som du har avlagt på finska eller svenska vid universitetet.
På museerna ordnas ofta också guidade rundvandringar på olika språk.
I tjänsten Uskonnot Suomessa (Religioner i Finland) finns information om religiösa samfund enligt ort.
Det syns överallt i den finländska kulturen, även i arbetslivet.
Importen är dock begränsad.
Rovaniemi stads invandrarbyrå
Du kan ansöka om studieplats i skolornas gemensamma ansökan på våren eller hösten.
När du besöker tjänstestället för att styrka din identitet ska du ta med dig ditt identitetsbevis och ansökningsbilagorna i original.
Flyktingrådgivningen ger asylsökande rättshjälp i asylprocessens första skede.
Rutterna för camping, paddling, vandring, cykling och övriga rutter i Karleby finns i karttjänsten på nätet.
Om man har flexibel arbetstid ska den anställda själv se till att han eller hon arbetar den tid som avtalats.
Om du behöver vård under samma dag ska du kontakta hälsostationen direkt på morgonen när den öppnar.
Efter moderskapsledigheten kan antingen modern eller fadern stanna hemma för att ta hand om barnet. Föräldraledigheten varar 158 vardagar.
Om föräldrarna har samma efternamn, blir detta även barnets efternamn.
har angett felaktiga uppgifter i medborgarskapsansökan eller medborgarskapsanmälan
Graviditeten avbryts med läkemedel eller med skrapning (kaavinta).
Om du har blivit utsatt för detta kan du få en öppningsoperation.
Det är viktigt att du känner väl till din bransch och de lagar som styr företagande.
Av speciellt vägande skäl kan abort göras även senare men då behöver du ett specialtillstånd från Valvira (Valvira).
Den andra föräldern får dock bestämma om vården och fostran av barnet när barnet är hos honom eller henne.
grammatik och vokabulär
Yrkeshögskolor, Universitet.
linkkiSettlementförbundet i Finland:
Finskt medborgarskap genom anmälan
Under den här tiden var Finland autonomt, vilket betyder att finländarna fick själva bestämma om många saker.
Då behöver du inte ett separat uppehållstillstånd för att arbeta.
Kontaktuppgifterna hittar på din kommuns hemsida.
Arbetskraftsbyråns informationstjänst för utbildning och yrkesval
Tillståndet måste sökas inom tre månader från barnets födelse.
Hjälp till offer för människohandel
Om du betalar för mycket skatt, får du skatteåterbäring.
Behandlingen på A-kliniken är konfidentiell.
Problem i äktenskapet?
Man ansöker om skilsmässa i tingsrätten.
Daghemmet är ändå inte en skola.
Ekonomi- och skuldrådgivarefinska _ svenska _ engelska
Att röra sig
Social- och krisjouren har öppet dygnet runt varje dag.
Detta innehåll finns inte på det språk som du har valt.
Fortsatt uppehållstillstånd för studerande
Laga inte mat om du är berusad.
Info om arbetskraftsutbildningfinska _ svenska
Klasslärarna i grundskolan, som undervisar årskurserna 1–6, har läst pedagogik.
En utredning över din försörjning i Finland
Tfn 029 56 61820
att få upplysningar om sitt hälsotillstånd, vårdens omfattning, riskfaktorer och alternativa behandlingsmetoder
De flesta finländarna är kristna.
Läs mer: linkkiJustitieministeriet:
Om översättningen görs av en auktoriserad översättare i Finland eller ett annat EU-land, behöver översättningen inte legaliseras.
Finländare går gärna rakt på sak i samtal.
Karens
Fastigheten utgörs vanligen av egnahemshuset och dess tomt.
Läs mer om detta på InfoFinlands sida När ett barn föds i Finland.
Man behöver alltså inte vänta tills betänketiden på sex månader har gått ut.
Handläggning av asylansökanfinska _ svenska _ engelska
Ring inte nödnumret vid vanliga sjukdomsfall.
En anställd vid arbets- och näringsbyrån gör den inledande kartläggningen
Moderskapsförpackningfinska _ svenska _ engelska
Om du inte kan betala räkningen på en gång, ska du kontakta inkassobyrån och komma överens om en betalningsplan för räkningen.
Övningar för allmänna språkexaminafinska
Ägarbostad
Rättshjälpsbyråerfinska _ svenska _ engelska
Ordna finansiering
I Varia ordnas även engelskspråkig undervisning samt finskspråkiga yrkesutbildningar särskilt avsedda för invandrare.
Omatila-tjänsten
Integrationsutbildning ordnas av kommuner, arbets- och näringsbyråer och många läroanstalter.
Din e-post används inte för några andra syften.
Ungdomar kan även söka bostad via ungdomsbostadsföreningen Rovaniemen nuorisoasunnot ry.
Barnets båda föräldrar är välkomna till rådgivningsbyrån.
När du flyttar utomlands för att bo där eller lämnar
Integrationsplanens längd beror på hur lång tid du behöver stöd för din integration.
en före detta finska medborgare
Polisen kan utfärda dig ett identitetskort för utlänningar om du har identifierats och din identitet har verifierats på ett tillförlitligt sätt.
Om du behöver hjälp med ett missbruksproblem (såsom alkohol- eller drogmissbruk), kan du kontakta din närmaste hälsostation.
Ibland kan också personer som inte omfattas av den finländska sjukförsäkringen ha rätt till ersättning från FPA.
Om föräldrarna utövar våld mot ett barn eller en ung, kan denne söka hjälp till exempel hos skolans hälsovårdare, vid familjerådgivningen eller FRK:s De ungas skyddshus.
Stöd för närståendevårdfinska _ svenska _ engelska
Ring 0295 000
Hälsovårdaren vid barnrådgivningen ger råd i frågor som rör små barns hälsa, uppväxt och utveckling.
Boka en tid hos preventivmedelsrådgivningens läkare eller hälsovårdare om du behöver preventivmedel (raskauden ehkäisy) eller om du överväger abort (abortti).
Yrkesutbildning för vuxna omfattar
Du kan samtidigt ansöka om medborgarskap för ett minderårigt barn som du har vårdnaden om.
Också den ungas föräldrar kan kontakta ungdomsstationen.
Du ska bifoga följande handlingar till din ansökan om uppehållstillstånd för studerande:
Finlands nationalmuseumfinska _ svenska _ engelska
Individens frihet syns starkt i den finländska lagstiftningen.
syskon eller halvsyskon
Målsättningen är att patienten kan återvända hem så fort som möjligt.
Ingen kultur eller religion får begränsa barns och ungas grundläggande rättigheter.
I Finland finns även vetenskapsbibliotek och läroanstalternas bibliotek samt olika slags specialbibliotek.
Finlands grundlag garanterar jämlikt bemötande för alla.
Preventivrådgivningfinska _ svenska
En brottsanmälan kan du göra på polisstationen.
Stadens hyresbostäder
linkkiFlyktingrådgivningen rf:
Seniorernas tjänster, serviceboendet och anstaltsvårdenfinska _ svenska
Om du flyttar till Finland tillfälligt har du vanligtvis inte rätt till den sociala tryggheten i Finland.
Öppettider och kontaktuppgifterfinska
Läs mer om högskoleutbildning på InfoFinlands sida: Högskoleutbildning.
Skilsmässan är officiell först när den andra ansökan har godkänts.
Du behöver också ett följebrev från kommunens socialväsen.
Om du inte blir antagen till integrationsutbildning på svenska kan du i vissa fall få stöd för frivilliga studier i svenska, om detta överenskommits i din integrations- eller sysselsättningsplan.
Studerande
Diskriminering och rasism
Du har rätt att jobba, fungera som företagare och studera i Finland.
Fölisöns friluftsmuseumfinska _ svenska _ engelska _ franska _ tyska
Förskoleundervisningfinska _ svenska
beväringar och civiltjänstgörare
Du kan fråga om detta på hälsostationen eller av skolhälsovårdaren.
Om du inte kan finska eller svenska kan du använda en tolk när du uträttar ärenden hos myndigheterna.
diplomingenjör
Allvarliga fall i samjour Uleåborgs universitetssjukhus (Oulun yliopistollinen sairaala OYS) kl. 21.00−8.00, tel. (08) 315 2655
Om du vistas i Finland i högst sex månader och din arbetsgivare är ett utländskt företag, behöver du i allmänhet inte betala skatt till Finland.
Daghem med vård på främmande språkfinska _ svenska _ engelska
Ditt röstningsställe har antecknats på meddelandekortet.
Rehabiliteringen genomförs på ett sätt som passar just dig.
Telefon: 040 8065 149
Mer information om ansökningsproceduren hittar du på InfoFinlands sida Fortsatt uppehållstillstånd.
Du kan också själv påverka vem din förmögenhet delas till.
Du kan själv söka information om lediga bostäder.
Arbetsavtalsmallar på olika språkfinska _ svenska _ engelska _ ryska _ estniska _ franska _ tyska
Barnets efternamn vid samboende
Arbetstagaren kan också be att orsaken till att anställningen upphört och en bedömning av arbetstagarens färdigheter och uppförande antecknas i intyget.
Samma person kan väljas till president högst två gånger.
Social- och krisjourenfinska _ svenska _ engelska
Karleby stadsbibliotek/huvudbiblioteket
Hyresvärden ansvarar till exempel för bostadens fasta inredning och ytmaterial.
I Finland värdesätts också demokrati och yttrandefrihet.
Specialsjukvård ges på centralsjukhus och universitetssjukhus.
I Vanda finns tjänster som är särskilt avsedda för äldre.
Personlig utvecklingsplan för kunnandet
Om du vill flytta till en familjemedlem som bor i Finland behöver du ett uppehållstillstånd.
Samtidigt är det bra att anmäla barnen till det nya daghemmet eller den nya skolan.
löneverifikat, d.v.s. ett lönebesked som arbetsgivaren gett.
Föräldradagpenningarna omfattar
Delaktighet
Museet för modern konst EMMAfinska _ svenska _ engelska _ ryska
Att ansöka om finskt medborgarskapfinska _ svenska _ engelska
När du känner igen grundläggande drag i den finländska företagskulturen kan du bättre betjäna dina kunder. Du har också bättre insikt i vad folk förväntar av dig.
Undervisningen på universitet är baserad på vetenskaplig forskning.
Adresserna är:
Om du flyttar utomlands för över sex månader anses din flytt vara permanent.
Också den tid som du har varit bosatt i något annat EU- eller EES-land kan delvis beaktas.
Avfall som inte får läggas i det egna husets sopbehållare kan föras till återvinningsstationer.
I grundskolorna ges även utbildning i finska som andraspråk (suomi toisena kielenä) till elever som har ett annat modersmål än finska, svenska eller samiska, och vars kunskaper i det finska språket inte är i nivå med modersmålet.
Fullmäktige väljs var fjärde år genom kommunalval (kunnallisvaalit).
Åklagaren överväger om hen väcker åtal.
Om du får avslag på din asylansökan eller ansökan om uppehållstillstånd har du rätt att överklaga beslutet.
I de flesta biblioteken finns en läsesal.
Återkallande av uppehållstillstånd
Fundera också på vilket kunnande du har fått från dina fritidsintressen eller andra erfarenheter.
När du är utomlands och har rätt till FPA:s förmåner ska du alltid anmäla ändringar i dina förhållanden till FPA.
Anmälningen ska göras till magistraten senast den 80:e dagen före valdagen.
Också handikapporganisationer tillhandahåller många slags hobbyverksamheter.
Dessutom ska ditt barn ha en finländsk personbeteckning.
Du kan ansöka om familjeåterförening även senare, men då tillämpas kravet på tillräcklig inkomst på er.
Undervisning för invandrare
utkomststöd
Målet är att alla, oavsett familjens inkomster, ska ha möjlighet att få en högklassig utbildning och växa till aktiva medborgare.
Vi följer användningen av sidorna, men samlar inte in några sådana uppgifter som kan kopplas till en person.
Förlossningssjukhusens jourmottagningfinska _ svenska _ engelska
Arbetsavtal
Helsingfors är Finlands huvudstad.
Förlovning
Mer information om rätten till hemkommun finns på InfoFinlands sida Hemkommun i Finland.
Om du vill studera vid ett vuxengymnasium ska du ta kontakt direkt med läroanstalten.
Den närmaste jourmottagningen för vuxna finns vid Jorv sjukhus.
Småbarns hälsa
I Finland tillämpas inga reservationsavgifter för bostäder.
Om du har ett tillfälligt uppehållstillstånd för arbete eller näringsidkande kan du ansöka om ett kontinuerligt uppehållstillstånd när du har vistats i Finland två år utan avbrott.
Vardagar kan tider till smärtjouren bokas enligt överenskommelse vid samtliga tandkliniker.
Busstidtabellerfinska _ svenska _ engelska
Mellersta Österbottens sommaruniversitetfinska
Du får göra ändringar i din bostad.
Dessutom kan du få vuxenutbildningsstöd (aikuiskoulutustuki).
På den här sidan finns allmän information om finländska seder.
På hälsostationerna finns läkarens, sjukskötarens och hälsovårdarens mottagningar.
Om du har barn och ska skilja dig, ta kontakt med barnatillsyningsmannen.
Språken i Infobanken är finska, svenska, engelska, ryska, estniska, franska, serbokroatiska, somaliska, spanska, turkiska, albanska, kinesiska, kurdiska (sorani), persiska och arabiska.
Karleby enhet
Ni
ditt barn som är under skolåldern är i privat dagvård; eller
linkkiInstitutet för hälsa och välfärd:
Tfn (09) 8306 220
Barn till en finsk medborgare
Du kan ringa TE-telefonservice då du behöver information om TE-byråns tjänster eller vägledning i tjänsterna på nätet.
Ungdomar och påverkan
tfn 040 0377 595
Finska undervisas som främmande språk och målet är en funktionell tvåspråkighet.
Barnet måste vara under 18 år gammalt och ogift den dag då beslutet om uppehållstillstånd fattas.
I huvudstadsregionen bor över en miljon människor.
Läs mer om ämnet: Registrering av uppehållsrätten för EU-medborgare.
Information om arbetarskyddfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
linkkiFritänkarförbundet r.f.:
Ofta innehåller de även anvisningar om användningen av gemensamma utrymmen i huset.
Läs mer på InfoFinlands sida Ingående av äktenskap i Finland, komihåglista och Äktenskapsförord.
Om det finns minst tre elever som befriats från religionsundervisningen och deras föräldrar kräver detta, ordnas undervisning i elevernas egen religion.
Vuxenutbildningscenterfinska
Om du har frågor kring stödtjänsterna för handikappade, kontakta handikappservicen vid Esbo stad.
Läs mer på InfoFinlands sida Barn vid skilsmässa.
Mer information om boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite får du av bland annat samkommunens servicestyrcentral, tfn 040 806 5093.
linkkiKanta:
Hemförsäkringar säljs av försäkringsbolag.
Du kan ansöka om uppehållskortet elektroniskt via tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Upphörandet av samboförhållandet kan påverka till exempel de stöd som FPA betalar och barnens dagvårdsavgifter.
Hjälp med att upprätta en affärsverksamhetsplan
Grundläggande utbildningfinska _ svenska _ engelska
du inte fyllt 18 år och inte har en vårdnadshavare i Finland.
Beslutsfattande och påverkan
Fråga på din studieort var du kan söka en studentbostad.
Tjänster för invandrarefinska _ svenska _ engelska
Inresetillstånd för utlänningarfinska _ svenska _ engelska
När du har ett möte ska du komma i tid.
Om ditt arbete pågår över tre månader ska du ansöka om ett säsongsarbetstillstånd hos Migrationsverket.
Anspråkslöshet
Om dina ekonomiska problem beror på spelproblem är det bäst att söka hjälp.
jobbsökningsförmåga och planerar sin framtid.
När du börjar på ett nytt jobb ska du lämna ditt skattekort till arbetsgivaren.
I vissa situationer kan studierna vid dessa läroanstalter dock vara kostnadsfria.
Om en brand uppstår, ring nödnumret 112.
Du har begått brott och du anses utgöra ett hot mot den allmänna ordningen och säkerheten.
Ring den kostnadsfria Jourhjälpen på tfn 116 117 innan du kommer till jourmottagningen.
Rådgivning och integration för invandrare
I Grankulla finns två gymnasier, ett finskspråkigt och ett svenskspråkigt.
Bostadsaktiebolagets ordningsregler anger när det ska vara tyst i huset.
Om aborten görs medicinskt doseras läkemedlet med 1–3 dagars mellanrum via slidan så att livmoderns börjar dras samman och töms.
Enligt finsk lag får ingen diskrimineras på grund av ett handikapp.
Tidsbeställningsnumret till tandvården i Helsingfors är (09) 310 51400.
Man kan till exempel komma överens om gemensamma regler med andra föräldrar.
Invandrarrådgivning
Svenska talas mest på Finlands väst- och sydkust.
Flerspråkiga ordböckerfinska _ svenska _ engelska
Om barnets vårdnadshavare är pensionerad kan han eller hon ansöka om en barnförhöjning på sin pension från Fpa.
Mer information om bouppteckningen får du från rättsväsendet och skatteförvaltningen.
Läs mer på InfoFinlands sida Den sociala tryggheten i Finland.
Detta betyder att man inte till exempel får slå eller lugga barn när de är olydiga.
Vid hindersprövningen utreder myndigheterna om det finns hinder för äktenskapet enligt Finlands lag.
Om du har ett Helmet-lånekort, kan du också låna böcker i Flerspråkiga biblioteket.
Karleby finns i Mellersta Österbotten invid Bottniska viken.
Studiehandledarna berättar om olika studiemetoder och om fortsatta studier.
Läs mer om barndagvård, förskoleundervisning och grundläggande utbildning på InfoFinlands sida Det finländska utbildningssystemet.
Invånarparker och klubbarfinska _ engelska
Lönen bestäms enligt kollektivavtalet.
du har tillräckliga kunskaper, färdigheter och resurser för den företagsverksamhet som du planerar
Grundläggande utbildning
Barnen studerar inte skolämnen och har inte lektioner.
Kravet på tillräcklig inkomst tillämpas dock inte på dig om ditt barn är en finsk medborgare.
Syftet med verksamheten är att stödja integrationen av invandrare, främja toleransen och acceptansen av mångfald, öka sysselsättningen, utveckla nya strategier och nätverka med aktörerna i regionen.
Om du vårdar ett barn som är yngre än tre år hemma kan du ansöka om hemvårdsstöd från Fpa. Skötaren kan till exempel vara barnets vårdnadshavare eller annan släkting.
Förteckning över yrkeshögskolorfinska _ svenska
Du hittar uppgifter om barns och ungas problem också på InfoFinlands sida Barns och ungas problem och Var hittar jag hjälp när barn eller unga har problem?
Omskärelse får inte göras utan smärtlindring som ges av läkare, och det ska göras i en steril miljö.
Registrerat parförhållande
I Finland gäller även en lag om likabehandling.
på skattebyrån
Det är föräldrarna som har ansvaret för att barnet går i skolan.
Om du har avlagt examen i Finland, behövs inte ett delbeslut av arbets- och näringsbyrån för ditt tillstånd.
Fyll i en ansökan och lägg till bilagorna.
Via dessa företag kan du även få en fast anställning.
Mångkulturell barndagvård i Rovaniemi betyder att alla barn beaktas likvärdigt och rättvist oavsett ålder, kön eller hudfärg.
Nylands arbets- och näringsbyrå hjälper invånare i Grankulla att söka jobb.
Skolhälsovårdaren tar hand om skolbarns hälsa.
Flyttkostnaderna beror på varifrån du flyttar och hur mycket saker du har.
Det finns 73 parkeringsautomater och du betalar parkeringsavgiften i en parkeringsautomat.
I bostadsrättsavtalet fastställs storleken på bostadsrättsavgiften, bruksvederlaget och övriga eventuella villkor.
Till exempel fysiskt våld eller stjälande är brott.
Finska medborgares rättigheter och skyldigheter
När du öppnar ett bankkonto har banken en lagstadgad skyldighet att fråga vad ditt konto ska användas till.
Mer information om FPA:s rehabiliteringar hittar du också på FPA:s webbplats.
Aktieägarens rösträtt, vinster och ansvar i företaget beror på hur många av bolagets aktier han eller hon äger.
Om du inte meddelar att du vill byta efternamn, behåller du ditt efternamn.
Grunden för näringslivet i Karleby är den internationella storindustrin.
Invandrarorganisationer
Mån–fre kl. 8.00–15.00; tis, ons, tors även kl. 17.00–19.30
För registreringen ska du lämna in ett legaliserat äktenskapsintyg i original till magistraten (maistraatti) i din hemkommun.
Om du är osäker på om smärtan är normal ska du fråga råd vid din egen rådgivningsbyrå.
Kontrollera att bostaden verkligen existerar, alltså att bostaden har samma adress som står på avtalet.
Dagverksamheten innefattar transport, en måltid, motion eller annan verksamhet.
De första 200 åren var staden en anspråkslös småstad.
Kommunerna i Finland kan vara antingen enspråkiga eller tvåspråkiga.
Klasslärarna i grundskolan, som undervisar årskurserna 1–6, har läst pedagogik.
Riksdagen
Arbets- och näringsbyråns arbetsplatssajtfinska _ svenska
I Finland finns också många föreningar som grundats av invandrare.
Mervärdesskatten (arvonlisävero) är en konsumtionsskatt som i Finland betalas för nästan alla varor och tjänster.
du har företagande som bisyssla och utvidgar företagsverksamheten till din huvudsyssla.
Men å andra sidan kan hyresvärden bestämma sig för att säga upp hyresavtalet, om han eller hon har en godtagbar anledning.
rådgivningen och kundtjänsten vid sektorn för fostran och utbildning:
Undervisnings- och kulturministeriet svarar för utvecklingen av och det internationella samarbetet inom utbildnings-, vetenskaps-, kultur-, motions- och ungdomspolitiken.
Läs mer: Skilsmässa.
I Esbo finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
Kontakta omedelbart fastighetsskötseln, disponenten eller hyresvärden.
Läs mer: Hyresbostad
Du har nytta av nätverk när du söker jobb.
Om du är medborgare i ett EU-land, EES-land, nordiskt land eller Schweiz och vill flytta till Finland för att starta ett företag, behöver du inget uppehållstillstånd.
Information om sexuellt likaberättigandefinska _ svenska _ engelska _ ryska
Detta kan exempelvis inkludera
I vissa fall kan du ändå få ett tillfälligt (B) uppehållstillstånd i Finland på grund av sällskapande.
Information för underhållsskyldigafinska
På utbildningsstyrelsens (Opetushallitus) webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
Enligt lagen om likabehandling måste arbetsgivare och utbildningsanordnare förbättra handikappade personers möjligheter att få arbete och utbildning.
+358 (0)29 497 152 (engelska)
När en närstående person avlider kan du få stöd och hjälp med din sorg vid hälsostationerna (terveysasema), på familjerådgivningen (perheneuvola), SOS-kriscentret för utlänningar inom Föreningen för mental hälsa i Finland (Suomen mielenterveysseuran ulkomaalaisten kriisipalvelu) samt hos församlingarna.
Flerfaldigt medborgarskap kan vara en fördel när man till exempel flyttar från ett land till ett annat.
tfn 016 322 2592
I stora städer finns också privata idrottsanläggningar.
Du kan också söka ersättning i efterhand med en blankett.
När du har avlagt yrkesinriktad grundexamen kan du söka dig till fortsatta studier antingen inom yrkesinriktad tilläggsutbildning, vid en yrkeshögskola eller vid ett universitet.
Arbetstagaren har rätt att få samma lön under semestern som under arbetet.
Information om privata hälsotjänster hittar du på sidorna Hälsa i Esbo och Hälsa i Helsingfors.
En familjemedlems död
Ett sådant utlåtande ger inte tjänstebehörighet i Finland, men det kan ändå vara till hjälp när man ansöker om ett arbete eller en studieplats, eftersom det beskriver innehållet i och nivån på utbildningen som man har avlagt utomlands.
Till musikskolorna ansöker man medelst inträdesprov en gång per år.
linkkiTuberkuloosi.fi:
VALMA-utbildningen kostar vanligen inget för den studerande.
Friluftsliv och vandringfinska _ svenska _ engelska
Modersmålsprovet kan skrivas i finska, svenska eller samiska.
Var och en har rätt att anmäla till polisen ett brott som ägt rum, alltså göra en brottsanmälan.
Uppehållstillstånd för arbetstagare är inte nödvändigt för alla arbetsuppgifter.
Hotell i Finlandfinska _ svenska _ engelska _ ryska _ kinesiska
Äktenskapet är alltid ett frivilligt val som ingen kan tvingas till.
Till apotekets tjänster hör också sidoapotek och apotekens tjänsteställen samt apotekets egen webbtjänst.
Mannen och kvinnan ansvarar båda för att ta hand om barnen och hemmet.
Besök fackevenemang i din bransch, gör frivilligarbete eller sök till ett mentorprogram.
anställa en arbetstagare
Preventivmedels- och familjeplaneringsrådgivningarna betjänar kvinnor och män i alla åldrar.
Du kan be om råd och hjälp också av Vailla vakinaista asuntoa ry.
Information om skidåkningfinska
Filmerfinska _ engelska
till en sund och trygg arbetsmiljö.
Det är vanligt att finländarna litar på andra människor och på myndigheter.
boendetjänster
Om du flyttar till en familjemedlem i Finland, krävs det ofta även att den person som bor i Finland har tillräckliga medel för att försörja sig själv och den familjemedlem som flyttar till Finland.
Läs mer på linkkiRovaniemi stad:
bostadsunderstöd i samband med militärunderstöd för värnpliktiga och civiltjänstgörare.
Samma person kan väljas till president för högst två mandatperioder efter varandra, det vill säga för tolv år.
Finska språket har sina rötter i de mellersta delarna av Ryssland, men har också inslag av baltiska och germanska språk.
Om du håller på att flytta till Finland, får du skattekortet från skattebyrån (verotoimisto).
Det betyder att det är bra att klä på sig åtminstone en täckjacka, ylletröja, mössa, handskar, halsduk och varma vinterskor.
På utrikesministeriets sida finns en lista över Finlands beskickningar utomlands.
För det behövs båda makarnas medgivande.
En anställning kan vara tidsbunden om orsaken är till exempel
Ta med dig pass, passfoto och originalexemplaren av ansökningsbilagorna.
Grundlagen
Läs mer på InfoFinlands sida: Efter grundskolan.
Finland tar som kvotflyktingar emot personer som har flyktingstatus enligt
Dra dig inte för att prata finska eller svenska med dina kollegor.
Ofta kan man få hjälp med att få barn.
Om du behöver särskilt stöd t.ex. på grund av handikapp ska du ansöka till utbildningen på våren, under ansökan till specialundervisning.
Studierna vid en yrkeshögskola (ammattikorkeakoulu) är praktiskt inriktade.
Förlossningssjukhusen i Helsingforsregionen är Kvinnokliniken (Helsingfors) och Jorv sjukhus (Esbo).
linkkiFöretagsfinland:
Då vårdas akuta sjukfall på jourmottagningen (päivystys).
Om du har ett tidsbestämt uppehållstillstånd med familjeband som grund kan det faktum att äktenskapet eller det registrerade parförhållandet upphör påverka uppehållstillståndet.
Hjälp i nödsituationer
Rådgivningstjänst för nordiska medborgarefinska _ engelska _ norska
Om du har avlagt en examen i Finland kan du få ett uppehållstillstånd för att söka arbete.
Verksamheten kan till exempel bestå av handledd motion, sång eller sysselsättning.
Om du väntar barn och känner att du inte klarar dig på egen hand kan du kontakta ett mödrahem (ensikoti).
Medborgarinstitut i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Det viktigaste redskapet för den som färdas på isen är isdubbar.
Läs mer: Gymnasium
Särdrag i undervisningen
Om du behöver psykoterapi som stöd för din arbets- eller studieförmåga, kan du eventuellt ansöka om rehabiliterande psykoterapi (kuntoutuspsykoterapia).
Om du redan befinner dig i Finland på någon annan grund kan du ha rätt att arbeta även om du inte har ansökt om ett uppehållstillstånd på grund av arbete.
Om du får uppehållstillstånd i Finland kan dina familjemedlemmar ansöka om tillstånd på grund av familjeband.
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) har du efter en självrisktid (omavastuuaika) rätt att söka sjukdagpenning (sairauspäiväraha) hos FPA (Kela).
Stöd för boendetfinska _ svenska _ engelska
Vid folkhögskolan kan man till exempel avlägga djurskötarexamen eller massörexamen.
Finansiering för ett företagfinska _ svenska _ engelska
Båda föräldrarna bär ansvaret för underhåll av ett barn under 18 år, även om de inte bor tillsammans.
Betala vattenavgiften till hyresvärdens eller husbolagets konto på samma gång som du betalar hyra.
Romppu
Barnbidraget betalas till den förälder hos vilken barnet bor officiellt.
Finlands Röda Kors kan inte bistå familjemedlemmarnas flygresor eller andra resor ekonomiskt.
I anslutning till folkhögskolan Työväen Akatemia i Grankulla finns en enhet för Humanistiska Yrkeshögskolan, där du kan avlägga yrkeshögskoleexamen för kulturproducenter.
Familjeplanering är helhetsbetonat främjande och upprätthållande av kvinnans och mannens sexuella hälsa.
Barnrådgivningens arbete omfattar hälsofrämjande arbete, förebyggande av sjukdomar och upptäckande av dem i ett tidigt skede samt uppföljning av och stöd för barnets helhetsbetonade psykiska, fysiska och sociala utveckling.
Servicepunkt
Information om arbets- och näringsbyråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Om du fallit offer för ett rasistiskt motiverat brott kan du göra en polisanmälan på nätet eller polisstationen.
I Helsingfors finns även många ungdomsgårdar, där de unga kan vistas på fritiden.
Försörjningsförutsättning för familjemedlemmar till personer som får internationellt skyddfinska _ svenska _ engelska
På den här sidan berättar vi om FPA:s stöd till studerande samt om penningunderstöd och stipendier.
I Finland finns ett rikt hobbyutbud för barn och unga.
De är avsedda för alla som vill lära sig att prata finska.
När du vill boka tid i tandvården ska du ringa tandvårdens tidsbeställning i din hemkommun.
Sambo med flykting
Innan du besöker magistraten kan du fylla i en registreringsanmälan som du kan ladda ned på adressen maistraatti.fi.
Flyktingen har förutsättningar att integreras i Finland.
Utbildningen är kostnadsfri för deltagarna.
Prövning av äktenskapshinder
Män som har fyllt 18 år har värnplikt (asevelvollisuus).
Ta med dig en identitetshandling och originalexemplaren av ansökningsbilagorna.
du har avlagt högskolestudier eller högskoleexamen utomlands.
Den finländska värdegrunden
_ lettiska
Om barnet har två vårdnadshavare, behövs varderas samtycke, i annat fall kan ingreppet inte göras.
Rehabiliteringsstöd är invaliditetspension på viss tid.
Regeringens verksamhetfinska _ svenska _ engelska
Att röra sig till sjöss
Frivilliga studier med stöd av arbetslöshetsförmånfinska _ svenska _ engelska
Finland anser att alla EU-länder är trygga för medborgarna.
Information om stöd- och serviceboendefinska _ svenska _ engelska
Du kan få rådgivning även om du inte är medlem i ett fackförbund.
Studeranden måste dock själv skaffa gymnasieböckerna.
Om barnet saknar tillräckliga färdigheter i finska eller svenska för att delta i undervisningen i klassen inleder han eller hon studierna i förberedande undervisning i en egen grupp eller i klassen enligt det egna studieprogrammet.
Den finska matkulturenengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ japanska _ italienska
Du kan avlägga examen för nöjaktiga eller goda språkkunskaper olika orter i Finland.
du har vistats två år utomlands utan avbrott.
På InfoFinlands sida Brott hittar du information om vad du kan göra om du blir utsatt för ett brott.
Ansök om en plats inom den kommunala småbarnspedagogiken från din egen kommun senast fyra månader innan du behöver den.
Som billigast kostar biljetten ungefär fem euro, som dyrast över tio euro.
Du kan också låta bostadsrätten gå i arv.
ditt barn provar på att återvända till skolan eller barnomsorgen.
Utlänningar som har rösträtt i kommunalval har även rätt att ställa upp som kandidat i kommunalval.
Barnet uppmuntras till självständigt tänkande.
Om barnets kunskaper i det finska språket inte är tillräckligt bra för studier i den finskspråkiga grundskolan, kan barnet få förberedande utbildning (valmistava opetus).
Domus Arctica-stiftelsens webbplatsfinska _ engelska
Tfn 116 117
Läs mer på InfoFinlands sida Utländska studerande i Finland.
Du kan få inkomstrelaterad dagpenning om du
Högskoleutbildning
Anonyma Alkoholister
Om du har avlagt examen i Finland kan du få ett tillfälligt uppehållstillstånd för att söka arbete.
Du ansöker om tillståndet vid Migrationsverkets servicesställen.
Om faderskapet erkänts före födelsen inleds behandlingen av faderskapsärendet först 30 dagar efter barnets födelse.
En full sopsäck ska tillslutas noggrant.
Läs mer på InfoFinlands sida Medborgare i nordiska länder.
I Helsingfors och Åbo finns en synagoga.
Sjukhusgatan 1
Om du har fått uppehållstillstånd på grund av behovet av skydd och får rätt till hemkommun i Finland, kan du utnyttja hälsovårdstjänsterna i din egen kommun.
Du kan fråga råd av hälsovårdaren (terveydenhoitaja) eller boka tid hos läkaren (lääkäri).
I registreringsblanketten finns en punkt där du kan be om att dina uppgifter registreras i befolkningsdatasystemet.
Om du vill hitta en arbetsplats i Finland ska du studera finska eller svenska.
Hur får jag arbetsintyget?
Läs mer: Äldre människors hälsa och Äldre människor.
Den snabba ekonomiska utvecklingen avtog i mitten av 1800-talet, men tog ny fart i slutet av århundradet tack vare industrialiseringen.
Ett friluftsmuseum kan till exempel vara en traditionell finländsk bondgård eller något annat område som gjorts om till ett museum.
Du kan ringa och boka tid.
I utlåtandet beskrivs examensnivån och innehåll samt för vilka uppgifter examen ger kvalifikationer i det land där du har avlagt examen.
På skattekortet anges en inkomstgräns och din skatteprocent beräknas utifrån den.
Tidsbeställning mån–fre 9–11
Få en födelseattest
Om du inte har rätt till de offentliga hälsovårdstjänsterna, kan du boka tid på en privat läkarstation.
Evenemangfinska _ engelska
Undervisning ges två timmar i veckan.
linkkiLapplands yrkeshögskola:
Hur grundar jag ett företag?
Om Migrationsverket ger dig ett positivt beslut på din asylansökan, får du uppehållstillstånd.
Läs mer på InfoFinlands sidor Stöd till gravida.
du har bott tillsammans med din sambo minst två år eller
Finnvera är ett finansieringsbolag som ägs av finska staten.
Det är bra att reservera minst en månad för att söka hyresbostad.
Om ni vill kan ni upprätta ett skriftligt avtal om umgängesarrangemanget.
linkkiFinnvera:
Anonyma Alkoholister (Anonyymit Alkoholistit) AA on är en kamratförening för män och kvinnor, där de delar med sig av sina erfarenheter av alkoholism och försöker hjälpa varandra att bli friska.
Det lönar sig att avsätta tid för bostadssökandet och undersöka olika alternativ.
Kurser i finska språket vid öppna universitetet
Fyll i ansökningsblanketten i Studieinfo.fi-tjänsten.
Bokbussarnas rutter och tidtabellerfinska
Make/maka till en flykting
Det betyder att barnet och familjen får stöd till exempel i skolan eller rådgivningen innan man kontaktar barnskyddet.
Om en person inte var medlem i kyrkan och inte ville ha en religiös begravning, förrättas en sådan inte.
Information om förskoleundervisningenfinska _ svenska
att skrämma, följa eller observera någon
Motionskarta över Karlebyfinska _ svenska
Vanligen börjar daghemsdagen på morgonen och tar slut på eftermiddagen.
Hälsostationerna når du genom att ringa till respektive hälsostations eget telefonnummer eller hälsorådgivningens telefonnummer (09) 839 10023 och väljer din hälsostation med hjälpa av knappsatsen.
Du kan hyra en bostad på den öppna marknaden.
Min granne klagar ständigt om oljud hos mig.
Kontrollera vilka kurser som är aktuella i institutets webbtjänst.
Din förälder eller mor- eller farförälder som är beroende av dig för sin försörjning
Om fördelningen av ägodelarna blir stridig, kan samborna i vissa fall ansöka om en bodelningsman hos tingsrätten som hjälper i bodelningen.
Om du vill kan du även skriva fler ämnen.
Ange om bearbetningar är gjorda.
Enligt lagen om jämställdhet ska myndigheter, arbetsgivare och läroanstalter främja jämställdheten mellan kvinnor och män.
Stödboendet hjälper dem att lära sig bo på egen hand och föra ett självständigt liv och stödjer dem i återhämtningen.
Utmätning betyder att myndigheten har rätt att ta en del av dina inkomster för betalning av skulder.
Juridisk rådgivning
Stadsfullmäktigefinska _ svenska _ engelska
Om du har avtalat om yrkesinriktad arbetskraftsutbildning i din sysselsättningsplan, kan du få förhöjd arbetslöshetsförmån.
Finland fick en egen lantdag 1906 och det första valet ordnades 1907.
Ring hälsostationen genast på morgonen för att boka tid.
Makarnas underhållsskyldighet
Information om registrering av fordonfinska _ svenska _ engelska
7 år
I staden finns dessutom två bokbussar som åker runt.
Du kan använda tolken när du själv önskar om du betalar kostnaderna och beställer tolken själv.
Jourmottagningen är öppen alla dagar dygnet runt
När vi lagar mat uppstår det mycket fukt i köket.
Personer som kommer till Finland som flyktingar kan ta del av integrationsrelaterade socialtjänster vid Rovaniemi stads invandrarbyrå.
Om du redan har avlagt en yrkesexamen eller en högskoleexamen, kan du inte söka till en yrkesutbildning i den gemensamma ansökan.
I Helsingfors finns flera begravningsplatser.
Myndighet
Vardagar kl. 15–08, fre–sön och helgdagar dygnet runt
I den privata sektorn krävs inget beslut om erkännande, men beslutet kan vara nyttigt då man söker jobb.
Även vuxna kan utbilda sig till ett nytt yrke eller komplettera sin kompetens.
Du ska bland annat registrera företaget, betala skatt och ordna bokföringen.
Om läkaren har skrivit ut ett elektroniskt recept (sähköinen resepti), kan du ta ut medicinerna på apoteket utan pappersrecept.
Fritid och hobbyer
I vissa skolor ges undervisningen på något annat språk än finska.
Finland var en del av Sverige i över 600 års tid från medeltiden till 1800-talets början.
Dessutom är de textade till finska och svenska.
Du kan få understöd för terapin ett år i taget under högst tre år.
Därefter kan eleven fortfarande läsa finska eller svenska som andraspråk, som S2-språk, om hen behöver stöd med språket.
I praktiken kan orsaken vara någon av följande:
Öva på att beskriva din bakgrund och din yrkeskunnighet med några meningar.
linkkiWebbtjänsten Suomi.fi:
Där kan du fråga om råd och få stöd i föräldraskapet och fostran av barn.
Civilvigsel förrättas i magistraten, religiös vigsel förrättas i en kyrka eller i något annat religiöst samfund.
Via Karleby löper riksväg 8 och 13.
Konstmuseetfinska _ svenska _ engelska
Bostadsrättsavtal
Det innebär att man på en stor lön betalar en större andel skatt än på en mindre lön.
Oberoende av vilket land du är medborgare i kan du i vissa fall arbeta i Finland utan uppehållstillstånd.
Om du arbetar och får lön eller är företagare behöver du ett finskt skattekort (verokortti).
En handikappad person bosatt i Karleby har rätt att erhålla de tjänster han eller hon behöver på samma grunder som de övriga invånarna i kommunen.
På sommaren ordnas avgiftsfri parkgympa på många håll i staden.
Boende i ägarbostad
Om du vill gå eller cykla i Vanda kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
Röstning
På biblioteket för synskadade Celia kan du låna ljudböcker, punktskriftsböcker, e-böcker och reliefbilder.
Om du ska gifta dig i Finland hittar du nyttig information på InfoFinlands sida Äktenskap.
inte under tiden har bott utomlands i över två år och
Innan du kan få körkort måste du delta i förarutbildning och avlägga förarexamen.
I Vanda ordnas LUVA-utbildning av Lumon lukio.
du är återflyttare, det vill säga återvänder till Finland från utlandet
I Vanda ges dagvård på finska, svenska, ryska och engelska.
Läs mer om den grundläggande utbildningen på InfoFinlands sida Grundläggande utbildning.
Om du är medborgare i ett EU-land, Liechtenstein eller Schweiz, behöver du inget uppehållstillstånd eller visum i Finland.
Du behöver bara visa upp ditt studentkort när du betalar för måltiden.
linkkiMuseiverket:
Fråga om mödrahemsverksamheten på din egen rådgivningsbyrå.
Teknik och trafik (ingenjör inom bilteknik, maskinmästare i sjöfartsbranschen)
Om du bor i höghus eller radhus, anmäl läckaget genast till journumret för husets servicebolag.
Ditt nummer sparas dock i en automat och du blir uppringd.
Registreringen av uppehållsrätten för en EU-medborgare och uppehållskortet för en familjemedlem till en EU-medborgare kan återkallas eller bli ogiltigt om:
När du startar ett eget företag kan du beviljas en startpeng som tryggar din utkomst under den tid då du inleder din företagsverksamhet.
Resor i Finland
Personer som har svårt att klara av de dagliga sysslorna utan hjälp, till exempel äldre eller personer med funktionsnedsättning, kan få ta del av hemvårdens stödtjänster.
Närmare information om ansökningstiderna hittar du via Studieinfo.fi-tjänsten.
Hjälp till invandrarkvinnor
I vissa situationer kan den förälder som bor med barnet ansöka om underhållsstöd (elatustuki) vid FPA.
Uppehållstillstånd för uppstartsföretagarefinska _ svenska _ engelska
linkkiSkatteförvaltningen:
Läs mer: Hälsa
Grundläggande informationfinska _ svenska _ engelska
Läs mer: Graviditet och förlossning.
På skattebyrån (verotoimisto) kan du sköta ärenden rörande skatter.
Abortfinska
moderskapspenning och särskild moderskapspenning
Utbildning som handleder för yrkesutbildning
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sortering av avfall.
Kontrollera vilket som är det vanligaste språket på din ort.
I Vanda finns flera museer.
Tillståndsbeslutet är avgiftsbelagt.
Ibland kan det vara artigt att nia.
Du kan ställa Migrationsverket (Maahanmuuttovirasto) en ansökan om att inte återkalla ditt uppehållstillstånd.
du lämnade felaktiga uppgifter när du ansökte om registreringen eller om uppehållskortet för en familjemedlem till en EU-medborgare
Mer information om Fennovoimas kärnkraftverksprojekt i Pyhäjoki:
Arbetsavtalet upprättas i två exemplar, ett till den anställda och ett till arbetsgivaren.
På ungdomsgården finns alltid någon vuxen, vanligen kommunens ungdomsarbetare eller ungdomsledare.
Därför är det viktigt att anmäla sig till kursen i god tid.
Polisen övervakar att trafikreglerna följs.
mån-tors kl. 8–15 och fre kl. 8–13
Arten av det arbete du ska utföra påverkar typen av tillstånd.
Reglerade yrkenfinska _ svenska _ engelska
Boka vigseltiden i magistraten eller tingsrätten i god tid för bröllopsdagen.
Vanda stad tillhandahåller olika tjänster för arbetslösa som hjälper dem att få kontakt med arbetslivet och hitta jobb.
Undervisning kan även fås på engelska.
På InfoFinlands sida Negativt beslut om uppehållstillstånd hittar du information om vad du kan göra om du får ett negativt beslut.
Centrumbiblioteket Oodi, adress: Tölöviksgatan 1
Du kan fråga råd i ärenden som rör utkomstskyddet för arbetslösa vid din egen TE-byrå.
linkkiAava:
Byråns tjänster är avgiftsfria.
Undervisnings- och kulturministeriet
Invandrarenheten
Språkkunskaper hjälper dig att förstå det nya samhället och underlättar skötseln av ärenden.
Du kan också förnya dina lån på Internet.
Gymnasier i Helsingforsfinska _ svenska _ engelska
Stöd och hjälp för kvinnor som utövar våld eller är oroliga för att de kommer att göra det.
Du har rätt att se bostaden i förväg och bostadsförmedlaren kan inte kräva att få betalt för detta.
Du kan få färdtjänst och följeslagare på resor som anknyter till arbete, studier eller fritid.
Familjer med främmande modersmål har vid behov rätt till tolktjänster.
I vissa kommuner har barnet rätt till 20 timmar småbarnspedagogik per vecka om den ena föräldern är hemma.
Du kan också välja att avlägga en engelskspråkig examen.
Av pappret görs dagstidningar eller wc-papper.
Det krävs även ämbetsbevis (virkatodistus), som du får från magistraten eller kyrkoherdeämbetet.
Operationen får inte göras om pojken motsätter sig.
grammatik och vokabulär
Boende i bostadsrättsbostad
Handläggning av ansökan är avgiftsbelagd.
Om du inte är van vid att använda en dator, fyll i en ansökan på papper och lämna in den på Migrationsverkets tjänsteställe.
Flyttsaker från EU-området
Gustav Vasa ville göra Helsingfors till en handelsstad som konkurrerar med Tallinn, och även holländska och tyska handelsmän flyttade till staden.
linkkiFinlands Psykologiförbund:
du är ett offer för människohandel och du inte har en hemkommun i Finland
TE-telefonservicefinska _ svenska _ engelska _ ryska
Om ditt barn insjuknar ska du kontakta hälsostationen vid behov.
I de största städerna kan det ta flera veckor eller månader innan man får en bostad.
Du kan ansöka om plats inom småbarnspedagogiken för ditt barn elektroniskt via tjänsten suomi.fi eller med en blankett på stadens webbplats (ansökan om småbarnspedagogik).
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, Skatteförvaltningen, FPA, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Sexuellt våld är
Dessutom ordnar även idrottsklubbar motion för små barn.
TE-byrån, FPA eller kommunen utreder din rätt till arbetslöshetstförmån eller utkomststöd under integrationsplanen.
Information om hemvårdsstödfinska _ svenska _ engelska
De som har fyllt 35 år kan söka sig till hälsocentralläkarens mottagning i sitt eget område.
Sambor kan dock upprätta ett testamente (testamentti) för det fall att någon avlider.
Företagsrådgivningfinska _ svenska _ engelska
Arbetsplatser i kommunernafinska _ svenska
etniskt ursprung,
Det är roligt och tryggt att röra sig i naturen när du väljer rutter som passar dig med hänsyn till din kondition och dina kunskaper och följer anvisningar.
Information om hälsorådgivningfinska
Finlands lagarfinska _ svenska _ engelska
Behandling av brottmål i Finland
Sambor har till exempel inte rätt att bo kvar i familjens gemensamma hem om det tillhör den döda sambon.
Information om Finland för utlänningarengelska
Om de övriga museerna hittar du information på Vanda stads webbplats.
Följande myndigheter hör till statens lokalförvaltning:
Socialhandledare 016-322 3123, 0400-695 037
Betjäning kan även fås via tolk på det egna modersmålet.
Utländsk examen i Finland
Också till exempel en släkting eller en bekant som har körkort och erfarenhet av att köra bil kan lära dig.
Anmäl dig som arbetslös arbetssökande
Via arbets- och näringsbyråerna kan man till exempel söka till kurser i det finska språket.
Ange också anställningens längd.
Avvisning och utvisningfinska _ svenska _ engelska
Juridiska tjänster är avgiftsbelagda men om du har små eller medelstora inkomster, kan du få helt eller delvis avgiftsfri rättshjälp från statens rättshjälpsbyrå.
Läs mer på InfoFinlands sida EU-medborgare och Nordisk medborgare.
Registerbeskrivning:
Varje avsnitt innehåller vokabulär- och grammatikövningar.
På slutet avlägger studerandena vanligtvis studentexamen.
Läs mer om hjälpmedel och tolktjänster på InfoFinlands sida Tjänster för handikappade.
Rovaniemi stads ungdomstjänster ordnar intressanta aktiviteter och intressant verksamhet för unga.
Utlandsfinländarnas intresseorganisationfinska _ svenska _ engelska
Fpa:s allmänna bostadsbidrag
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta tjänsten Omatila (Omatila).
På hälsostationen bedöms din situation.
Parktanten övervakar och leder barnen som leker i parken.
Man ansöker till förberedande undervisning för gymnasiet under sommaren på webbsidan Opintopolku.fi.
I Finland är en person man sällskapar med inte en familjemedlem enligt lagen.
Läs mer om att söka jobb i Finland på sidan Var hittar jag jobb?
Information om papperslöshetfinska _ engelska _ franska _ arabiska
Studier
I regel har alla finska medborgare som fyllt 18 år rätt att rösta vid val.
Verksamheten sker på finska.
du har känt till det innan köpet.
Evenemang och festivalerfinska _ engelska
I Finland föder kvinnorna oftast på sjukhus.
tfn (09) 8393 5534
Under prövotiden kan arbetstagaren bedöma om arbetet lämpar sig för honom eller henne och arbetsgivaren kan bedöma om arbetstagaren är lämplig för arbetet.
Om du vill ansöka om finskt medborgarskap måste du kunna finska, svenska eller i det finska teckenspråket.
Information om finländska sederengelska _ spanska _ kinesiska _ tyska _ portugisiska
Om en person dör utanför sjukhuset ska du genast anmäla ärendet till polisen eller en läkare.
Besök på Nupoli är kostnadsfria och konfidentiella.
Vad gör jag när en vattenkran läcker?
Läs mer om den inledande kartläggningen och integrationsplanen på InfoFinlands webbplats Integration i Finland
Högskolorfinska _ engelska
År 1950 hade Esbo 25 000 invånare och 15 år senare redan 65 000 invånare.
Till exempel kan barnets lärare kontakta barnskyddsmyndigheterna.
Ett barn får finskt medborgarskap också om hen föds i Finland och inte får medborgarskap i något annan land av sina föräldrar.
E-post kan du skicka till adressen: kirjaamo.lappi(at)te-toimisto.fi
Att människor behandlas på olika sätt innebär inte alltid att det är fråga om diskriminering.
Du kan få betjäning på finska och engelska.
Det är vanligtvis det tryggaste sättet.
Filmer på främmande språk har vanligen finsk- och svenskspråkig textning.
Öva på att besvara allmänna frågor som ingår i en anställningsintervju.
Befolkningen är framför allt koncentrerad till de stora städerna och tätorterna.
Läkaren skriver en remiss till undersökningar på barnlöshetspolikliniken.
I Finland har polisen ansvaret för att reda ut brott och lämna dem till åtalsprövning.
Den allra ljusaste månaden är juni.
Mer information om barnets rättigheter i olika åldrar finns på InfoFinlands sida Barns och ungdomars rättigheter och skyldigheter.
För en vistelse som varar ett år ska du alltså ha 6 720 euro i disponibla medel.
Utan tillstånd får du inte göra några ändringar, även om du skulle bekosta renoveringen själv.
Denna summa är vanligen några procent av bostadens pris.
Många organisationer erbjuder även utbildning, rådgivning och olika stödtjänster.
Barn till en utländsk medborgare
I Finland finns det fem ansvarsområden för arbetarskydd som lyder under Regionförvaltningsverket (RFV).
om du är under 17 eller över 40 år gammal
Delta och påverkafinska
Ett sådant får du på biblioteket.
Upplevelser som kan orsaka ett trauma är exempelvis:
I nödfall kan du använda kommunala tjänster även om Esbo inte är din hemkommun.
åldringar
Finland är indelat i kommuner.
Om du kommer klockan 12.10 är du försenad.
Du har brutit mot inresereglerna och din ansökan har avslagits, till exempel på grund av skenäktenskap.
Asuntosäätiö har delägarbostäder i Esbo.
i familjedagvård eller
Via programmet kan du få en mentor, som stödjer dig i sökningen efter arbete eller utbildningsplats eller i att starta eget företag.
Finland var på den tiden en del av Sverige.
SERI-stödcentret
Du kan uppskatta din skatteprocent med Skatteförvaltningens skatteräknare.
Nämn också om du är rädd för att din närstående kommer att skada sig själv.
Alla som ansöker om en förskoleplats ska lämna in en ansökan om förskoleundervisning.
Vi hoppas att få se känslofyllda, intelligenta, smarta och roliga videoklipp.
Det är ändå inte alltid möjligt att få en plats på en annan skola.
Penningsummans storlek beror på vilket land du återvänder till.
Asylsökande har vanligtvis inte tillgång till offentlig hälsoåvård exempelvis på hälsocentraler.
blir utsatt för hot, eller om en närstående till dig blir utsatt för hot
Utnyttja sociala medier i jobbsökningen
Välj efternamnet tillsammans med din make eller maka redan när ni ansöker om prövning av hinder mot äktenskap.
På bankernas webbsidor finns det låneräknare.
linkkiHRM:
Läkaren bedömer din synskada och därefter kan du få hjälpmedel i form av medicinsk rehabilitering.
Om ett barn under 10 år insjuknar akut kan barnets mamma eller pappa stanna hemma för att ta hand om barnet.
Hejdå.
Även om arbetstagaren har sådan utbildning som krävs för yrket redan när anställningen inleds, uppmuntrar många arbetsgivare sina anställda att skaffa sig mer utbildning.
du har flyttat till Finland
Planera företagets finansiering noga innan du grundar företaget.
Du kan få behovsprövad rehabilitering om hälso- och sjukvården konstaterar att du har en skada eller sjukdom som kräver rehabilitering.
Telefon
Skillnaderna i olika skolors studieresultat är små och nästan alla avlägger grundskolan inom den utsatta tiden.
du får det allmänna bostadsbidraget
Du kan byta ut ditt körkort till ett finskt körkort på Ajovarmas serviceställen.
Läs mer på InfoFinlands sida Uppehållstillstånd för make eller maka.
information om arbetsplatser i Europafinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ norska
Läs mer: Att grunda ett företag
Meddela bostadsaktiebolaget eller disponenten, i praktiken vanligtvis allra först fastighetsskötseln, om det finns ett sådant fel i din bostad vars åtgärdande åligger bostadsaktiebolaget.
Stadsstyrelsen representerar kommunen: den använder stadens yttranderätt och vidtar olika juridiska åtgärder för staden.
Information om jämlikhet och likabehandling hittar du på InfoFinlands sida Jämställdhet och jämlikhet.
Berätta om mobbning för läraren eller rektorn.
Naturbruk- och miljöområdet
Arbete kan ge dig partiell rätt till social trygghet i Finland.
Yrkesutbildning ges av yrkesläroanstalter (ammatillinen oppilaitos), specialyrkesläroanstalter (erityisammattioppilaitos) och av vuxenläroanstalter (aikuisopisto).
Din rätt till bostadsbidrag och utkomststöd kan du få reda på hos FPA.
Telefonnumret till TE-telefonservice är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
Många museer har fritt inträde på den internationella museidagen 18.5.
Kom ihåg att anmäla dig också direkt efter studier, arbetskraftsutbildning eller en period med sysselsättningsstöd.
Tidsbeställningen till tandkliniken vid Grankulla hälsostation mån–fre:
FPA kan även ordna rehabilitering som behovsprövad rehabilitering (harkinnanvarainen kuntoutus).
Om samboförhållandet upphör på grund av att den ena parten dör, ärver samborna inte varandra.
tel. 06 826 4111
För uppgifter inom den offentliga sektorn (kommun eller stat) krävs ofta examen på en viss nivå, till exempel en högre högskoleexamen.
Om familjens yngsta barn är under tre år, kan barnets förälder få hemvårdsstöd (kotihoidon tuki) när han eller hon vårdar barnet i hemmet.
Mer information om gymnasieskolorna och den förberedande undervisningen för gymnasiet fås av stadens undervisningstjänster.
Grundläggande utbildning och gymnasiumfinska _ svenska _ engelska
Om du har hemkommun (kotikunta) i Finland kan du utnyttja de offentliga tandvårdstjänsterna.
När du har en hemkommun har du rätt att använda denna kommuns tjänster såsom till exempel offentliga hälsovårdstjänster.
EU-länderfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
Om du måste sköta ärenden med myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du använda en tolktjänst.
I Helsingfors finns ett svenskspråkigt universitet och en svenskspråkig yrkeshögskola.
Förvärvsinkomsten beskattas progressivt, d.v.s. ju större inkomster man har, desto mer skatt betalar man.
På full arbetslöshetsförmån ställs även andra villkor.
I Grankulla ordnas kurser i finska och svenska av Grankulla medborgarinstitut.
Arbetspension utomlands
Köparen har rätt att läsa köpebrevet före dagen då köpet genomförs.
Museer och traditionsarbetefinska _ svenska _ engelska
Företagets skatter betalas på basis av de beskattningsbara inkomsterna, vars belopp man uppskattar på förhand.
Missbruksproblem
Yrkesutbildning Högskolor
Lochteå tandklinik
Tfn: 09 31013300
+358 (0)29 497 150 (finska)
Det finns även vissa andra fall där du kan ansöka om skilsmässa enligt Finlands lag.
Läs mer: Missbruksproblem.
I början av CV:t kan du tillfoga en sammanfattning eller profil där du beskriver din bakgrund och din kärnkompetens med några ord.
Studielånet är ett lån som finska staten ger garanti för åt studeranden.
När du arbetar i Finland måste du betala skatter.
Grankullavägen 7
Om du jobbar inom byggbranschen behöver du också ett skattenummer (veronumero).
Det är viktigt att hålla sina löften och tala sanning.
Du kan skicka in ansökan till tingsrättens kansli per post eller via e-post.
På julen sjunger man julsånger och umgås med familjen och andra nära och kära.
Läs mer: Mental hälsa.
Pensionen kan utbetalas till vilket land som helst.
På sidan finns även information om att bo i hyresbostad och om sådant som rör flytten.
Hyresboende
De ger också yrkesvägledning.
att tvinga någon att tigga eller begå brott
Diskutera på finska
Att beställa ett arbetspensionsutdragfinska _ svenska _ engelska _ ryska _ estniska
Grundläggande information
Brottsofferjouren (RIKU) har till uppgift att främja brottsoffrets ställning samt ställningen för deras närstående och brottsmålsvittnen.
utbildning
InfoFinland-tjänsten ger dock ingen rådgivning och du kan inte ringa InfoFinland.
Tfn (09) 839 22133
I vissa fall kan banken även kräva andra utredningar av identiteten, om du har en notering i din handling som anger att din identitet inte har kunnat fastställas.
Där finns böcker på fler än 60 olika språk.
Också många sjukskötare har rätt att skriva ut vissa läkemedel.
Mer information får du på Migrationsverkets (Maahanmuuttovirasto) webbplats.
Förlossning
Läs mer under rubriken Stöd för frivillig återresa.
Utkomstskydd för arbetslösafinska _ svenska _ engelska
I grundskolan studerar barnen många obligatoriska ämnen.
Det finns också andra alternativ än ägarbostad och hyresbostad.
Skogarna, kärren, ängarna, åkrarna, älvarna och de små insjöarna skapar en bild av Lappland och Rovaniemi, vars uttryck och stämning ändras och förnyas i takt med årstiderna.
I Helsingfors finns många museer.
Ett registrerat partnerskap kan ändras till äktenskap vid magistraten.
Invånarhus Kylämajafinska
Dessa dagar kan inte överföras till modern.
Information om skatteförvaltningenfinska _ svenska _ engelska
Skyldighet att delta i landets försvar eller bistå i det.
Ungdomsgården är centret för ungdomsarbetet i respektive område.
Vid hälsostationerna vårdas även könssjukdomar (sukupuolitauti).
Nästan alla begravningsplatser i Finland ägs av evangelisk-lutherska församlingar men man kan få en gravplats även om man inte är medlem i den evangelisk-lutherska kyrkan.
Handel bedrevs längs med Bottniska vikens kust och jordbruk, jakt, fiske och sälfångst var även viktiga näringar.
Johan Ludvig Runeberg (1804–1877) är en viktig finländsk skald.
Till exempel sjukskötare kan avlägga högre yrkeshögskoleexamen inom rehabilitering.
Flickor kan få stöd och råd i Flickornas hus (Tyttöjen talo) och pojkar i Pojkarnas hus (Poikien talo).
Om du har blivit utsatt för könsstympning kan du få en öppningsoperation.
Du måste alltså ännu betala hyra för juli.
De lär sig också att respektera andra människors språk och kulturer.
Antalet ledamöter beror på invånarantalet i valkretsen.
Rättigheter
Fastighetsförmedlare och privatpersoner annonserar bostäder som de säljer i lokaltidningar (såsom Lapin Kansa) och på Internet.
Du kan hämta ditt bibliotekskort vid vilket HelMet-bibliotek som helst.
Folkhögskolorna ordnar mycket undervisning för invandrare.
Familjemedlemmar och andra anhöriga kan vara:
På språkcaféerna talar vi finska, så det är bra om du redan kan lite finska.
Då kan du söka till utbildningen i den kontinuerliga ansökan.
Museer och utställningarfinska _ svenska _ engelska
linkkiPatent- och registerstryrelsen:
linkkiFöretagsFinland:
Registrering av utlänningar 029 55 36 300
De är till exempel familjer som bildas av två kvinnor eller två män samt familjer med fler än två föräldrar
Karleby är en gammal sjöstad som erbjuder mångsidiga möjligheter för utfärder och friluftsliv.
ett heltidsarbete under de tider då ingen undervisning ordnas vid läroanstalten, vanligen under sommar- och vinterlov.
Lapplands yrkesinstitut
Många företag erbjuder förmånliga utlandsprefix.
Om ditt hem har fler än en våning måste du räkna ytan separat för varje våning.
Den internationella mötesplatsen Trapesa erbjuder rådgivningstjänster.
Familjerådgivningens telefonnummer: 044 730 7640.
Personligt resekort kan du köpa vid serviceställena.
Folk i Finland är aktiva motionärer och olika motionshobbyer kan hjälpa dig att bli bekant med människor och få nya vänner.
Fadern är vanligtvis med på förlossningen. Stödpersonen kan också vara en släkting eller en vän.
De finns i hus som ägs av ett bostadsaktiebolag.
Hemtjänsterna är hjälp med vardagssysslor, till exempel med att tvätta sig, klä på sig och måltider.
Naturhistoriska centralmuseetfinska _ svenska _ engelska _ ryska
Du ska inte heller ringa nödnumret om du vill fråga polisen (poliisi) till exempel om ett tillståndsärende.
Om du behöver hjälp eller stöd i mental- och/eller missbruksfrågor, boka tid till en psykiatriskötare.
du har begått två eller flera brott
Du hittar skilsmässoansökan på tjänsten suomi.fi.
Du kan få handledning i jobbsökningen.
Mitt hem i ett höghus(pdf, 6,56 MB)finska _ engelska _ ryska _ somaliska _ arabiska
Klubbarna räcker vanligen ett par timmar.
Finskans grammatikfinska _ svenska _ engelska _ ryska _ spanska _ tyska _ japanska
När du har hittat ett jobb kan du ansöka om uppehållstillstånd.
När du ska sköta ärenden vid polisens tillståndsenhet, kan du boka tid på förhand på polisens webbplats.
Komihåglista för nya studerande
Verksamheten i lekparkerna är avgiftsfri och öppen för alla.
Helsingfors tingsrättfinska _ svenska _ engelska
Ryssland erövrade Finlands område från Sverige 1808–1809.
Information om bibliotekets öppettider och tjänster finns på dess webbplats.
Om du är medborgare i något annat land behöver du ett uppehållstillstånd för studier.
FöretagsFinland ger dig information om olika finansieringsalternativ.
Vissa yrkesläroanstalter och gymnasieskolor ordnar förberedande utbildning före studierna.
I vissa fall kan du få folkpension även innan du fyllt 65 år.
Presidenten väljs i presidentval.
Läs mer: Grundläggande utbildning.
I tjänsten Enter Finland kan du betala med nätbankskoderna för en finsk bank eller med kreditkort.
Förskoleundervisningen ges av lärare med utbildning i pedagogik i minst 700 timmar om året, dvs. cirka fyra timmar om dagen, enligt skolans arbetstider.
Anställningsvillkoren bestäms enligt arbetslagstiftningen och kollektivavtalet.
Om du redan är försäkrad i ett annat land, behöver du ett intyg A1/E101 över försäkringen.
Du kan också göra brottsanmälan på internet om brottet i fråga är ringa och du inte behöver omedelbar hjälp av polisen.
Ibland hittar man ingen medicinsk orsak till den.
om din vistelse i Finland är tillfällig, beroende på hur länge vistelsen varar.
Fritid
Att söka uppehållstillstånd på grund av familjebandfinska _ svenska _ engelska
Detta beror på hurdant och hur långt arbetsavtal du har samt från vilket land du har kommit till Finland.
Läs mer: När du väntar barn.
Vid yrkesskolorna finns många olika områden som du kan studera.
När du öppnar ett bankkonto behöver du ett pass, ett identitetskort för utlänningar eller någon annan officiell identitetshandling.
Boende, arbete och försäkring
Nödnumret 112 fungerar i alla EU-länder.
Kalkkers håller öppet kl. kl. 22–6.
Miehen linja (Miehen linja) hjälper invandrarmän som har problem med våld.
Skattedeklaration och beskattningsbeslutfinska _ svenska _ engelska
Hem och familjfinska _ svenska _ engelska _ ryska _ estniska
Samtidigt hade man emellertid även kontakter med handelscentra i öst och den ortodoxa kyrkan.
Sjukvårdskortet ska vara giltigt under hela din vistelse i Finland.
Tfn 09 816 42439
A-klinikens tjänster är avsedda för personer som har fyllt 25 år.
Under den yrkesinriktade arbetskraftsutbildningen får du samma förmån som när du är arbetslös.
Trafiklänkar
På sidan Städer hittar du kommunerna som finns i InfoFinland på en karta.
Läroplikten upphör i slutet av det läsår då barnet fyller 17.
Teater och danskonst i Karlebyfinska _ svenska _ engelska
pensioner
Det beviljas även för dem som köper eller bygger ett egnahemshus.
Du behöver inget Apostille-intyg om du har en allmän handling som utfärdats av en myndighet i ett EU-land.
tfn (09) 816 33333
För handikappade och personer som återhämtar sig från mentala problem erbjuds bostäder som beaktar invånarnas särskilda behov.
Du får ingen ersättning för läkemedel som du köper utan recept.
Du kan också vara vårdledig på deltid.
Barn och unga serveras mat i daghem och skolor.
När man har beslutat något tillsammans förväntar sig både de anställda och arbetsgivaren att alla gör det man kommit överens om.
Tjänsten omfattar inte arbets- och näringsbyråns kurser.
Sortera avfallet enligt material.
Du får handledning och råd om att ansöka om socialtjänster och förmåner avsedda för handikappade samt med att fylla i blanketter.
Om situationen kräver det har du rätt att besöka hälsostationen inom tre vardagar efter att du kontaktade hälsostationen.
I den här listan har vi samlat de vanligaste ärendena som du måste ta hand om när du har kommit till Finland.
Projektet Sport för alla (Sporttia kaikille-hanke) ordnar idrottsklubbar, turneringar och läger för barn och ungdomar med invandrarbakgrund.
Vaccinering av personer över 65 år utförs vid seniorrådgivning.
linkkiVåldtäktskriscentralen Tukinainen:
Tillstånd till att avbryta graviditetenfinska _ svenska
Barns rättigheter
Settlementföreningen Rovalan Setlementti ry/MoniNet
På Miehen Linja kan du prata på finska, svenska, engelska, franska och grekiska eller medelst en tolk på ditt modersmål.
I ett samboförhållande behåller vardera part sin egen egendom.
Läs mer på InfoFinlands sidor Fackförbund och Arbetslöshetsförsäkring.
Romppu är settlementföreningen Rovalan Setlementti ry:s drog- och rusmedelsmottagning för ungdomar i Lappland.
Där kan man även studera finska och andra språk.
Familjen till ett barn som är under ett år gammalt kallas till barnrådgivningen minst nio gånger.
du har avtalat om utbildningen i din sysselsättningsplan med arbets- och näringsbyrån.
Missbrukarvårdfinska _ engelska
Läs mer: Förlossning.
I Finland tillhandahålls högskoleutbildning av yrkeshögskolor och universitet.
Kontaktuppgifter finns på webbplatsen för Helsingfors stad.
Ortodoxa kyrkan i Finland är landets näst största religiösa samfund.
Du kan också ha studier som hobby.
Många religiösa samfund är verksamma i Esbo och Helsingfors.
Tillfälligt boende.
Kommunerna har beskattningsrätt, det vill säga rätt att uppbära kommunalskatt av sina invånare.
Om du emellertid börjar arbeta i ett annat land eller reser utomlands för över ett år, kan din rätt till den sociala tryggheten i Finland upphöra.
I Esbo ordnas språkkurser i finska och svenska av Esbo arbetarinstitut, Esbo vuxengymnasium, Luksia och Axxell.
Valet av kvotflyktingar påverkas till exempel av följande faktorer:
Ledd motion
du inte har råd att skaffa en ägarbostad på samma område.
I Helsingfors finns en engelskspråkig Al-Anon-grupp.
Barnskyddet stöder familjer i problematiska situationer
om du har en förälder som är finsk medborgare,
Utländska studerande kan ansöka om olika penningunderstöd för finländska högskolor.
Fråga mer om omskärelse på rådgivningsbyrån, en hälsostationsläkare, skolhälsovårdaren eller skolläkaren.
skådespelare
Om du får en studentbostad kan du vanligen bo i den under hela studietiden.
Fadern får vårdnad om barnet om föräldrarna ingår ett avtal om gemensam vårdnad och faderskapet har erkänts.
Framskridandet av en HIV-infektion kan bromsas med läkemedel.
När du pratar med någon, ta ögonkontakt med personen du pratar med.
linkkitvguido.com:
Gör en ansökan innan ditt föregående uppehållstillstånd går ut.
Närings-, trafik- och miljöcentralerna (NTM-centralerna)
Typiska lönetillägg i Finland är erfarenhetstillägg, övertidstillägg och skiftarbetstillägg.
linkkiArbets- och näringsministeriet:
Du kan söka till en yrkeshögskola då du har avlagt en yrkesskola, gymnasiet eller studentexamen i Finland eller i ett annat land.
Högskolorfinska
Lapplands öppna universitetfinska _ engelska
Om du blir bostadslös, ta då kontakt med servicestället för socialarbete på ditt område.
Information om att bo i delägarbostadfinska _ svenska _ engelska
Om din bostad har skadats, till exempel till följd av brand eller vattenskada, kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Efternamnet påverkas inte av att samboförhållandet eventuellt upphör.
Om du har ett tillfälligt uppehållstillstånd på grund av familjeband kan du ansöka om ett kontinuerligt uppehållstillstånd när en familjemedlem till dig ansöker om ett kontinuerligt uppehållstillstånd.
Sveaborgfinska _ svenska _ engelska
Hälsostationerna enligt stadsdelfinska _ svenska _ engelska
Du kan på förhand fråga myndigheten om detta.
utsänd arbetstagare.
Läs mer om efternamn vid skilsmässa på sidan Skilsmässa.
Ledd motion ordnas till exempel av olika idrottssällskap som ofta drivs med frivilligarbete.
De har tystnadsplikt. De berättar inte om dina saker för andra myndigheter.
Operationen görs på sjukhus och återhämtningen tar vanligtvis 1–2 dagar.
tfn 020 634 0200
Om du är medborgare i något annat land har du med ditt uppehållstillstånd för studerande rätt att arbeta i begränsad omfattning, om arbetet är
Till förskoleundervisningen anmäler man sig via Esbo stads webbplats.
Om du är medborgare i ett nordiskt land behöver du inte uppehållstillstånd i Finland.
Du behöver uppehållstillstånd för arbetstagare om du arbetar till exempel som:
På hösten är det också mörkt, eftersom solen går ner tidigare än på sommaren.
Guiden God hyressed(pdf, 546 kB)finska _ svenska _ engelska
Karleby evangelisk-lutherska församlingssammanslutnings invandrararbete stöder invandrares integrering i det finländska samhället.
När allt finns på papper kan både den anställda och arbetsgivaren kontrollera i avtalet vad man gemensamt har avtalat.
Hjälp och information för personer som drabbats av etnisk diskrimineringfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska
Telefonnumret till Global Clinic i Helsingfors är 044 977 4547.
Kontaktuppgifterna till närmaste socialbyrå hittar du på din hemkommuns webbplats.
Av redogörelsen ska det åtminstone framgå
11 procent har något annat modersmål.
Det är viktigt att man regelbundet följer Wilma.
Nationella audiovisuella arkivet visar nya och gamla filmer från hela världen.
Dessutom finns det några tvåspråkiga universitet där du kan läsa på svenska.
Du inte lämnar landet frivilligt inom den tidsfrist som meddelats för dig.
linkkiMellersta Österbottens Familjerådgivningscentral:
Lagen förbjuder även diskriminering på grund av könsidentitet eller uttryck för kön.
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Om du har sökt asyl eller vistats i något annat EU-land (eller i Schweiz, Norge, Island eller Liechtenstein) innan du kom till Finland, behandlas din ansökan inte i Finland.
Mer information hittar du på Vanda stads webbplats.
Jourmottagningen är avsedd för situationer där man behöver omedelbar vård.
Fråga om ansökningstiderna vid medborgarinstitutets eller arbetarinstitutets studiebyrå.
I detta fall fastställer Migrationsverket barnets medborgarskap.
Invånarhuset Kivenkolo
Jämställande av nivån på en högskolexamenfinska _ svenska _ engelska
Höghuslägenheter och radhuslägenheter är bostadsaktier.
Underuthyrning
Du har lättare att sköta dina ärenden med myndigheter, följa nyheter, få nya bekantskaper och vänner.
Lokgränden 7
Läs avtalet noga innan du undertecknar det.
Finlands officiella språk är finska och svenska.
EU-medborgare som är i det finska rösträttsregistret kan också ställa upp som kandidat i Finlands Europaparlamentsval.
I hjärtat av staden, i det anrika Rooska gården, finns K.H.Renlunds museum.
Duschen, vattenkranarna och toalettstolen hör alltid till utrustningen.
Du hittar kontaktuppgifterna på Väestöliittos webbplats.
Tjänster för barnfamiljer
Ansökan om uppehållstillstånd för specialist
Studiestöd till utländska studerandefinska _ svenska _ engelska
Anställningsrådgivning för invandrarefinska _ svenska _ engelska
Finland som stöder företag bedömer ditt företags affärsmodell, kunnande och förmåga att få verksamheten att växa.
Om du insjuknar akut eller råkar ut för en olycka och inte kan vänta tills hälsostationen öppnar, kontakta jourmottagningen.
att de utländska studierna tillgodoräknas som en del av en finländsk examen.
När du är gravid
Fråga din arbetsgivare hurdana språkkunskapskrav som gäller på den arbetsplats som du vill söka.
Den sexuella skyddsåldersgränsen för barn är 16 år.
Kontaktuppgifterna finns under länkarna nedan.
På MoniNets webbplats finns länkar till olika webbsidor där du kan studera finska på egen hand.
Till befolkningen i Finland hör olika slags minoriteter som till exempel har ett annat modersmål, en annan kultur eller religion än majoriteten av finländarna.
Flickornas husfinska
Hushållsavfall
Konfessionslös begravningsplatsfinska
Fråga mer hos FPA:s center för internationella ärenden.
Om äktenskapet inte ingås inom denna tid måste hindersprövningen göras på nytt.
Med undersökningarna utreds varför en graviditet inte har börjat.
På viktiga bemärkelsedagar (födelsedagar, äktenskap, pensionering) uppmärksammar arbetskamraterna och arbetsgivaren festföremålet med en liten present eller en blombukett.
Du kan begära att FPA utreder din rätt till de offentliga hälsovårdstjänsterna.
I Vanda anordnas samtalsklubbar på finska också på Silkesportens verksamhetscenter (Silkinportin toimintakeskus) och Kafnettis och Myyrinkis boendeträffpunkter (Kafnetin ja Myyringin asukastila).
När barnet börjar i dagvården fyller man tillsammans med familjen i blanketten Uppgifter om invandrarbarn.
Priserna för den privata småbarnspedagogiken varierar.
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
Varken staden eller andra hyresvärdar är skyldiga att erbjuda dig en bostad.
Begränsningarna beror på vilken sorts läkemedel det är fråga om och från vilket land du tar med dig läkemedlet till Finland.
Språkkunskaper och finskt medborgarskapfinska _ svenska _ engelska
Detta kallas för Dublinprocessen.
Integration av invandrarefinska _ svenska _ engelska
Vid dem kan man inte avlägga yrkesinriktade studier.
Läs mer: Fritidsverksamhet för barn och unga.
om ni har bott tillsammans minst fem år.
Du kan skriva på finska, svenska eller engelska.
I den förberedande undervisningen ges undervisning i finska och i grundskolans ämnen.
När Finland blev självständigt år 1917 blev Helsingfors huvudstad i republiken Finland.
Kontrollera om dina nuvarande försäkringar, som hemförsäkringen, är tillräckliga även för den nya bostaden.
När du fyllt i ansökningen, kom ihåg att följa ditt konto i Enter Finland-tjänsten.
Säkerhetslås skyddar mot inbrottstjuvar
Det är dock inte givet att man får asyl, utan varje fall utreds separat.
I yrkeshögskolor kan du studera inom många områden.
Invandrare har rätt till en inledande kartläggning.
Förlängning av visum i Finland
I många bibliotek hittar du böcker på engelska, tyska, franska, italienska, spanska, estniska och ryska.
InfoFinland utvecklas i samarbete med finansiärerna.
Om du upptäcker att din hörsel blivit sämre, boka en tid för en hörselundersökning på hälsostationen i ditt område eller hos en privatläkare.
När du flyttar till Finland bedömer FPA alltid först om din flytt till Finland är stadigvarande boende i den mening som avses i lagarna om social trygghet.
En anställd får inte särbehandlas i arbetslivet på grund av graviditet eller föräldraskap.
Mottagning /Lochteå
Du kan få permanent uppehållstillstånd (pysyvä oleskelulupa) (P), om
Lapplands landskapsbibliotek/alla verksamhetsställen linkkiLapplands landskapsbibliotek/alla verksamhetsställen:
Om någon i din familj utövar våld mot dig eller hotar dig med våld, kan du kontakta ett skyddshem.
Moderskaps- och föräldrapenning kan betalas till exempel till mödrar som mitt under föräldrapenningsperioden flyttar till ett annat EU/EES-land eller Schweiz för mindre än ett år.
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus i Esbo och på Barnkliniken i Helsingfors.
Sponsringslöften eller kontoutdrag från privatpersoner, såsom släktingar, bekanta eller arbetsgivare, godkänns inte.
Om den ena föräldern har ensam vårdnad om barnet, kan den föräldern ensam bestämma vilket trossamfund barnet ska höra till.
Faderskapet fastställs av magistratet.
Läs mer:
Familjerådgivningfinska _ svenska _ engelska
Tfn (09) 816 35900
Uppehållstillstånd för företagare
Frivilligarbete kan dessutom bli en bra hobby.
På biblioteken i Helsingfors ordnas språkkaféer, där man kan öva sig i att prata finska.
Om din sambo har uppehållstillstånd i Finland och bor i Finland kan du få uppehållstillstånd i Finland på grund av familjeband.
människor som återhämtar sig från problem med den mentala hälsan och missbrukarproblem.
På InfoFinlands sida Bostadsbidrag finns information om det bostadsbidrag som FPA betalar.
ett hyresavtal som gäller tillsvidare eller
Utkomststöd söks hos FPA.
Du kan söka till en högre YH-examen på ett främmande språk med en separat ansökan.
Några museer, som till exempel Helsingfors stadsmuseum, har alltid fritt inträde.
Dessa finns till exempel på arbetarinstitut, bildkonstskolor, musikskolor och kommunernas ungdomsväsende.
linkkiTrasek ry.:
Därför bor många finländare i ganska små bostäder.
att vägra vård
Om du är rädd inför förlossningen, prata om det på rådgivningsbyrån.
Uppsägningstiden börjar i allmänhet först från slutet av den månad då avtalet sägs upp.
Läroavtalsutbildning ges till exempel vid många vuxenutbildningscentra (aikuiskoulutuskeskus).
Ekonomin och bokföringen ska granskas i slutet av perioden.
I Vanda finns två yrkeshögskolor (ammattikorkeakoulu), Laurea och Metropolia.
I Helsingfors är bostäderna i allmänhet dyra, men priserna varierar mycket mellan olika områden.
Ofta hjälper det redan att tala om dessa saker med familjen eller vänner. Ibland behövs det även annan hjälp.
Kristelefon för arabisktalande: 09 2525 0113.
Ta kontakt med polisen på din hemort.
Böckerna är ofta dyra.
Grundskolan är vanligen nioårig: skolan börjar i årskurs 1 och slutar i årskurs 9.
Ohjaamofinska _ svenska _ engelska
Alla som köper varor och tjänster är konsumenter.
Tillräcklig finansiering och noggrann planering är nödvändiga.
Dem kan du fråga om råd och få stöd i föräldraskapet och fostran av barn.
Med myndigheter avses till exempel polisen, FPA, arbets- och näringsbyrån eller tjänstemän vid Esbo stad.
16 år
Vuxengymnasietfinska
Lågstadiet omfattar årskurserna 1–6, högstadiet årskurserna 7–9.
I den andra valomgången kandiderar de två kandidater som fick flest röster vid första valomgången.
Bifogat till beslutet finns en anvisning om hur du överklagar.
linkkiJämställdhetsombudsmannens byrå:
För fiske krävs fiskelov, med undantag för mete och pilkning.
Om du är EU-medborgare behöver du inte uppehållstillstånd i Finland.
Serviceguide för seniorer(pdf, 1 MB)finska
Du kan köpa ett graviditetstest på apoteket.
Oy
Om du är kund vid arbets- och näringsbyrån kan du fråga om språkkurser i finska och svenska vid arbets- och näringsbyrån.
Ansökningstiden är vanligtvis i januari.
I Helsingfors finns även svenskspråkiga teatrar.
Valmansföreningen ska ha minst tio medlemmar.
Läs mer: Kulturer och religioner i Finland.
Du kan styrka din identitet vid Migrationsverkets tjänsteställe eller utomlands vid Finlands beskickning.
Om du för in en bil från ett land utanför EES-området behöver du också ett förflyttningstillstånd innan du kan använda bilen.
vardagen känns tung
Största delen av undervisningen på högskolorna ges på finska.
Människor framhäver sig inte i gruppen; de talar inte högljutt och skryter inte.
på nätet
minst en av föräldrarna arbetar i Finland och därmed omfattas av den sociala tryggheten i Finland.
Finlands flyktinghjälp r.f. är en organisation som strävar efter att främja de grundläggande rättigheterna för flyktingar.
Elektronisk ansökningsblankett för dagvårdenfinska _ svenska _ engelska
arbetspraktik.
Om du av någon anledning inte till exempel lyckas få en läkartid utanför arbetstiden, ska du komma överens med din chef om att du är borta och hur du ersätter din frånvaro.
I den öppna ansökan ska du berätta vad du kan och hurdana uppgifter du skulle kunna utföra.
Mer information om hälsovården i Finland får du på InfoFinlands sida Hälsa.
Om du blir arbetslös ska du anmäla dig hos TE-byrån senast den första dagen av din arbetslöshet.
De anställda ska också själva sörja för arbetssäkerheten.
I vissa höghus finns det också en brandsläckare i trappuppgången.
Global Clinic bedriver verksamhet i följande städer:
Huruvida du får lön under familjeledigheten beror på ditt kollektivavtal.
Permanent uppehållsrätt för EU-medborgare ansöks separat från Migrationsverket.
Jämfört med många andra länder har arbetstagare i Finland långa semestrar.
På magistraten kan du, under förutsättning att villkoren för detta uppfylls, även få en finsk personbeteckning, om du inte redan fick en sådan då du beviljades uppehållstillstånd eller din uppehållsrätt för EU-medborgare registrerades.
Läs mer på InfoFinlands sida Utkomstskydd för arbetslösa.
Privata hyresbostäderfinska _ svenska
I integrationsplanen antecknas åtgärder som främjar din integration.
Staten stöder boende i ägarbostad genom att gå i borgen för privatpersoners bostadslån.
Rovaniemi har alltid haft rollen som porten till Lappland och staden har varit det administrativa centret för Lapplands län ända sedan år 1938.
Europass är ett allmäneuropeiskt CV, alltså en allmäneuropeisk meritförteckning.
När du flyttar till Finland på grund av familjeband, har du obegränsad rätt att arbeta och studera i Finland.
År 1640 flyttades Helsingfors till stadens nuvarande plats på Estnäs.
Staden Rovaniemi är belägen mellan två stora älvar, Ounasälv och Kemi älv, och har blivit ett framstegsvänligt och internationellt centrum för handel, administration och utbildning.
Man kan även träna sina finskakunskaper i invånarlokalen i Kivenkolo.
Du kan få yrkesinriktad rehabilitering om du har sådana hälsoproblem som hindrar dig från att arbeta.
Utbildningsområden i yrkesutbildningenfinska _ svenska
Reglerade yrken och ansvariga myndigheterfinska _ svenska _ engelska
någon annan högskoleexamen
Hälsostationen och centralsjukhuset bekostar de hjälpmedel som ges som medicinsk rehabilitering (lääkinnällinen kuntoutus).
linkkiRättsväsendet:
Med läkaren eller psykologen kan du samtala konfidentiellt. De har tystnadsplikt.
Den humanistiska och pedagogiska branschen (teckenspråkstolk)
När du flyttar ska du meddela din nya adress till biblioteket.
Läs mer om VALMA-utbildningen på InfoFinlands sida Utbildning som handleder för yrkesutbildning.
Diskrimineringsombudsmannen och diskriminerings- och jämställdhetsnämnden övervakar att människor inte diskrimineras på grund av sitt etniska ursprung.
Föreningen Monika-Naiset Liitto har en jourtelefon för invandrarkvinnor som blivit utsatta för våld.
Du får mer information om stöd för närståendevård vid socialbyrån på din egen ort.
registreringsintyg över uppehållsrätten (oleskeluoikeuden rekisteröintitodistus) (om du är medborgare i ett EU-land)
Ta med dig identitetsbevis om du ska köpa personligt resekort.
Information om den förberedande utbildningen får du vid rådgivningen och kundtjänsten vid Stadin ammatti- ja aikuisopisto.
eventuella reparationsarbeten
Fråga mer hos FPA.
När du ingår ett hyresavtal i Finland, ska du nästan alltid betala en hyresgaranti.
Välfärds- och servicepunkten Olkkarifinska
Läs mer: Finlands förvaltning, Val och röstning i Finland
Vanda tillhör samkommunen Helsingforsregionens trafik (HRT) (Helsingin seudun liikenne -kuntayhtymä (HSL)), som ordnar kollektivtrafiken i huvudstadsregionen.
Vid NewCo Helsinki får du råd och hjälp med att starta ett företag.
Skolhälsovårdaren har hand om skolbarns hälsa.
Vissa delägarbostäder byggs med statligt stöd.
Om du vill fortsätta dina studier i Finland kan de studier som du avlagt utomlands tillgodoräknas med hjälp av akademiskt erkännande.
I detta fall kan du ansöka om visum i detta lands beskickning.
Om du, av anledningar som du inte själv kan påverka, inte hinner ansöka om uppehållstillstånd inom tre månader, kan du ändå ansöka om familjeåterförening.
Kurserna i svenska hittar du genom att klicka på länken på tjänstens startsida.
Om du måste låta utföra ändringsarbeten i din bostad eller montera fasta hjälpmedel i bostaden kan du få ersättning för dessa av kommunen.
Museer och slottfinska _ svenska _ engelska
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Sambo till en utländsk medborgarefinska _ svenska _ engelska
Sexuell hälsa och prevention
På den här sidan finns information om den bosättningsbaserade sociala tryggheten som hör till FPA:s ansvarsområde.
Ring inte nödnumret om det inte är en nödsituation.
I Finland finns flera organisationer som arbetar för att förbättra handikappade personers ställning i samhället.
På Helsingfors stads webbplats finns mer information om var du kan köpa fisketillstånd.
Du kan till exempel få ett brandlarm avsett för hörselskadade och en texttelefon för att kunna bo tryggt i ditt hem.
Startpeng (starttiraha)
I gymnasiet tas inga terminsavgifter ut.
Du kan också boka tid hos barnrådgivningens (lastenneuvola) psykolog eller en läkare på din egen hälsostation.
I vissa fall kan frivilligarbete vara en del av din integrationsplan.
Medlaren är oftast en anställd vid socialbyrån, barnrådgivningen eller familjerådgivningen.
föräldrarnas gemensamma efternamn eller
Temperaturen kan t.ex. dagtid vara -10 Celsiusgrader och ibland till och med -20 grader.
Läs mer: Skilsmässa.
Vi läser tillsammans för kvinnor
Avgifter i egnahemshus
Skattenummerfinska _ svenska _ engelska
Vad gör tolken?
Läs mer om dessa och andra viktiga frågor som en företagare bör veta på InfoFinlands sida Företagarens skyldigheter.
Det kan hjälpa att tala med en hälsovårdare (terveydenhoitaja), läkare (lääkäri) eller en psykoterapeut (psykoterapeutti).
Dessa är Sveaborg, Gamla Raumo, Petäjävesi gamla kyrka, Verla träsliperi och pappfabrik, Sammallahdenmäki fornlämningsområde, Struves kedja och Kvarkens skärgård.
Vid problem i äktenskap eller parförhållande får du hjälp av Mellersta Österbottens familjerådgivningscentral som underhålls av Karleby kyrkliga samfällighets och Mellersta Österbottens social- och hälsovårdssamkommun Soites familjerådgivning.
Studentbostäder
Vid akuta krissituationer inom familjen kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys), som har öppet dygnet runt varje dag.
Vem kan ingå äktenskap?
Den här sidan är avsedd för dig som är medborgare i något annat land är ett EU-land, Norge, Island, Schweiz eller Liechtenstein.
Om det görs av icke-medicinska orsaker, inkräktar man på en pojkes fysiska integritet.
Om du vill att ditt barn ska börja i svenskspråkig dagvård, förskola eller skola, fråga om möjligheterna i din hemkommun.
Om du är EU-medborgare eller nordisk medborgare:
yrkesexamina
I vissa städer finns en poliklinik för könssjukdomar där könssjukdomar behandlas.
Läs mer: Hyresbostad
I krissituationer får man även hjälp vid Vanda stads social- och krisjour (sosiaali- ja kriisipäivystys), som har öppet dygnet runt.
Mer information om hur du gör medborgarskapsanmälan hittar du på Migrationsverkets webbplats.
Du kan också betala kursavgiften på Internet om du har webbankkoder till Handelsbanken, Sparbanken Optia, Nordea, Andelsbanken eller Danske Bank.
Rådgivningsbyråernas tidsbokning och rådgivning
Diskrimineringsombudsmannen
linkkiKiasma:
Om inkomstgränsen överskrids ska du beställa ett nytt skattekort.
Läs mer: Gymnasium.
Kontakta rådgivningsbyrån när du upptäcker att du är gravid.
Ungdomscentralen (Nuorisoasiainkeskus) erbjuder många idrottsmöjligheter till 9–18-åriga barn och unga.
Klubbarna för att lära sig tala finska är avgiftsfria.
Ta med dig dina arbetslöshetsförmånerfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
Om du vill fördjupa dina yrkeskunskaper kan du avlägga högre yrkeshögskoleexamen (ylempi ammattikorkeakoulututkinto).
Universitet och institutioner har olika ansökningstider.
Mån.–fre. kl. 9–15
Du behöver vanligtvis inte skicka in dina arbetsintyg i förväg till arbetsgivaren, men det är bra att ta med dem till anställningsintervjun för det fall att arbetsgivaren vill se dem.
I Grankulla finns en evangelisk-luthersk kyrka med två församlingar, en finskspråkig och en svenskspråkig.
Läroavtal (oppisopimus) innebär inlärning i arbetet.
Rehabilitering för arbete
Notera att utländska handlingar måste vara legaliserade för att man utgående från dem ska kunna föra in personuppgifter i befolkningsdatasystemet.
När du har en arbetsplats ska du kontakta läroavtalsbyrån (oppisopimustoimisto) i din region.
Du kan skicka in din fråga via webblanketten på finska, svenska eller engelska.
Man kan inte ansöka om att bli kvotflykting via myndigheterna i Finland.
Övriga avgifter
Tidsbokning vardagar kl. 12–13
Hälsovårdaren på barnrådgivningsbyrån ger råd i frågor som gäller små barns hälsa, tillväxt och utveckling.
Restiden med tåg till Helsingfors är cirka fyra timmar.
Du kan i regel komma till jourmottagningen genom att först kontakta jouren via telefon.
Välj ansökningsblankett utifrån grunden för din ansökan om nytt tillstånd.
Även ett barn som föds i Finland behöver ett uppehållstillstånd i Finland.
Flyktingen utgör inget hot för Finlands säkerhet.
Tiondeklasserna i Vanda finns i östra och västra Vanda vid Varias verksamhetsställen och vid Lumo gymnasium (Lumon lukio).
Barnets mor är finsk medborgare.
Yrkesinriktad rehabiliteringfinska _ svenska _ engelska
Allemansrätten ger inte rätt att skräpa ner i naturen, skada träd eller växter, störa eller skada fågelbon eller fågelungar, köra motorfordon utan markägarens tillstånd eller bygga ens tillfälliga byggen.
I Vanda finns två kulturhus: konserthuset Martinus och allaktivitetscentret Myrbackahuset.
Du kan anmäla dig till vårens kurser i början av året och till höstens kurser i slutet av sommaren.
Boende i ägarbostad
Du kan vara partiellt vårdledig tills barnet har gått ut årskurs två.
Däremot följs inlärningsresultaten upp med urvalsbaserade bedömningar.
Varje hälsostation har ett eget telefonnummer för tidsbokning, som man kan ringa för att boka tid till sjukskötare eller läkare.
Om din granne ofta och på ett allvarligt sätt bryter mot ordningsreglerna, kan du kontakta disponenten eller hyresvärden.
I Finland kan du få personbeteckningen även vid magistraten eller skattebyrån på din hemort.
Läs mer om Fpa på InfoFinlands sida Viktiga myndigheter.
Föräldrar som har gemensam vårdnad beslutar tillsammans om många saker. Dessa är barnets
Då anger lagstiftningen till exempel hur lång hyrestiden i bostaden är och hur man kan avstå från bostaden.
service och reparationer
uppdrag som sakkunnig
På Apotekareförbundets (Apteekkariliitto) webbplats kan du söka information om apoteken på din hemort och deras öppettider.
som har rösträtt i kommunalval,
Sådana är till exempel boendetjänster, arbetsverksamhet och dagverksamhet.
linkkiPatent- och registerstyrelsen:
Diskriminerings- och jämställdhetsnämnden
Det lönar sig att ansluta sig till en arbetslöshetskassa, eftersom den inkomstrelaterade dagpenningen är större än det vanliga utkomstskyddet för arbetslösa.
Om du vill flytta till Finland behöver du vanligtvis ett uppehållstillstånd.
Sveaborg och Stora Räntan är också historiska sevärdheter.
Vid behov kallas du till undersökning.
Finland tillhör Schengenområdet.
Allmän information om boende:
Om faderskapet inte fastställs är barnet officiellt faderlöst och då ansvarar modern ensam för underhåll och vård av barnet, även om ni bor tillsammans.
Sådan praxis är dock ovanlig på arbetsplatser.
linkkiExpatFinland:
Kontrollera uppgifterna i skattedeklarationen.
är 16–67 år
Du kan skriva till Väestöliittos mångkulturella kunskapscenter på dari, kurdiska (sorani), persiska, finska, ryska, engelska eller svenska.
Du kan ansöka om besöksförbud hos polisen eller i tingsrätten (käräjäoikeus).
Gymnasierna och gymnasiernas hemsidorfinska
Sådana betalningar är till exempel skatter, hälscentralsavgifter och dagvårdsavgifter.
FPA betalar in studiepenningen på ditt konto månatligen.
Ta med ett ID-kort och ditt uppehållstillstånd.
minst tre års arbetserfarenhet från samma område som din examen och du har inhämtat din arbetserfarenhet efter att du har avlagt examen.
Läs mer om hjälpmedel för synskadade och hörselskadade på InfoFinlands sida Handikappade personer.
Finlands grannländer är Ryssland (i öster), Norge (i norr), Sverige (i väster) och Estland (i söder).
Hur stort stöd du får beror på hur mycket hjälp du behöver.
Specialyrkesexamen (erityisammattitutkinto)
Vid tidsbeställningen bedöms även om du behöver vård av läkare eller hälsovårdare.
Kompetenscenterfinska
Kontaktuppgifter till utbildningsväsendetfinska _ engelska
Läs mer: Äldre människor.
En utredning över företagsverksamheten (om du är egenföretagare)
Handikappade
Lekparks- och eftermiddagsverksamhet för skolbarnfinska _ engelska _ ryska _ somaliska _ arabiska
Läs mer: Brott.
Handikappade barns skolgång
Om det inte finns några medicinska skäl till omskärelsen kan den inte utföras inom den offentliga hälsovården.
Finskt medborgarskap är inte samma sak som uppehållstillstånd.
Man badar bastu med såväl familjemedlemmar och vänner som med affärspartner.
Du kan tala finska, svenska eller engelska.
På vintern ska man klä sig varmt i Finland.
Skeppsvarv fanns bland annat i Kaustarviken, Svartskär och Soldatskär.
Läs mer på InfoFinlands sida Till Finland för att arbeta.
Missbrukararbete
Du kan också boka tid hos en privat gynekolog. Privatläkares tjänster är avsevärt dyrare för kunden.
trettondagen 6.1
arbets- och näringsbyråerna,
Om en anställd till exempel vill hålla en bönestund under arbetsdagen ska detta göras under de avtalade pauserna.
Det är viktigt att du har ett arbetsintyg från alla anställningar i Finland.
Kontaktuppgifter:
I Finland betraktas som familjemedlemmar
Peluuri är en hjälptelefon för personer med spelproblem, deras närstående och andra som möter spelproblem.
I ordningsreglerna anges vanligtvis till exempel tiderna för när det ska vara tyst i huset.
Du kan få hjälp på flera olika språk.
Historiafinska _ svenska
Du behöver inte boka tid på jourmottagningen.
ett tidsbestämt hyresavtal.
Telefon: (06) 8287 701
Att rösta i kommunalvalet är ett viktigt sätt att påverka.
Du kan söka invalidpension hos FPA.
Om du är sjuk en lång tid ska du ta reda på om rehabilitering kan vara till nytta för dig.
Förlovningen är ett löfte om äktenskap.
linkkiArbetsministeriet:
Vissa dagar är allmänna lediga dagar i Finland.
Hjälp för ungafinska _ svenska _ engelska
Du får vård även vid en långvarig sjukdom.
Om du har ett företag i Vanda, kan du bli medlem i Vanda Företagare.
Med familjeledighet avses
Köparen kan betala handpenningen åt säljaren i det skedet då köpet förbereds.
På InfoFinlands sida Avfallshantering och återvinning hittar du information om sopsortering.
Servicestället i Rovaniemi
För att skydda kunderna uppges inte klinikens adress eller öppettider offentligt.
Äldre människor kan anlita tjänster som tillhandahålls av vanliga hälsostationer.
KOSEKs experter hjälper bland annat med att utarbeta en affärsverksamhetsplan och att ansöka startpeng.
Närmare information hittar du på hälsostationernas egna webbplatser.
Arbets- och näringsministeriet
På Vanda stadsbibliotek anordnas språkcaféer (kielikahvila), där man kan öva på att prata finska.
Målet är att med hjälp av motion förbättra både den psykiska hälsan och den fysiska konditionen.
Läs mer: Teater och film.
Makarna kan även ansöka om ett helt nytt efternamn som deras gemensamma namn.
Detta betyder att en 16-åring är försäkrad mot ålderdom, arbetslöshet och arbetsoförmåga och att sjukförsäkringsersättningen betalas till den unga själv, inte dennes föräldrar.
Självständighetens tidiga år 1917–1945
missbrukarvård
Du får mer information på InfoFinlands sida under rubriken Hälsovårdstjänster i Finland.
Presidenten är Finlands statsöverhuvud.
I Finland har en arbetstagare rätt:
Även Marthaförbundet och Finlands flyktinghjälp erbjuder bostadsrådgivning åt invandrare.
Utred bostadens skick och andra frågor
Fuktproblem
Läs mer: Sexuell hälsa och prevention.
Tfn (09) 816 52044 och (09) 816 52043
Biblioteken har böcker och annat material på flera olika språk.
Ansökan är fritt formulerad men datum, underskrift och dina personuppgifter ska finnas med.
Gör anmälan till handelsregistret och skattemyndigheten
Hur länge användarna stannar kvar på sidorna
Karleby mödra- och skyddshemfinska
Tfn (09) 816 5800
Lagarna stiftas av riksdagen.
De kan dessutom tillhandahålla andra tjänster.
Du kan ta reda på om det är möjligt att registrera en hemkommun i Finland för dig vid magistraten på din hemort.
Vem sköter företagarnas intressebevakning i Finland?
Psykiatriskötarna har mottagning på hälsostationerna.
Skidåkning
I Finland har program på främmande språk text på finska eller svenska, med andra ord kan man också titta på dem på originalspråket (oftast engelska).
Om arbetet är uppenbart farligt kan den anställda vägra att utföra det.
Bostadsrättsbostad
De hjälper dig att utveckla affärsidén och planera affärsverksamheten.
Adress
På läkemedelsförpackningen står det sista användningsdatumet.
Caisafinska _ svenska _ engelska
Du ansöker till yrkesinriktad arbetskraftsutbildning antingen i arbets- och näringsbyrån eller med en elektronisk blankett på internet.
(Eurooppalainen viitekehys EVK) Denna skala omfattar följande nivåer:
En familj kan ha barn eller bestå av ett barnlöst par.
Följande kan få allmänt bostadsbidrag
Om du har arbetat i andra länder som Finland inte har ett socialskyddsavtal med, måste du själv ta reda på om du har rätt att få pension från dessa länder.
Din försörjning behöver inte vara tryggad i följande fall:
Undervisning i finska för barn
Mer information hittar du på HNS webbplats.
Fråga mer om senioruniversitetet i kansliet för närmaste öppna universitet.
På vintern är det ofta halt ute.
Östra Nylands rättshjälpsbyrå (Itä-Uudenmaan oikeusaputoimisto) betjänar invånarna i Vanda.
Du kan avlägga en yrkesinriktad grundexamen antingen
Manslinjen
FPA:s bidrag är avsedda för personer som omfattas av Den sociala tryggheten i Finland.
Fråga mer på FPA.
Information om arbetarskydd och råd vid problemfinska _ svenska _ engelska
Finland är en republik.
Ansökan om skilsmässa görs i två skeden.
C2 – ASE 6
Öppningsoperationen kan även göras i mitten av graviditeten.
Innan du anmäler dig till examen ska du göra dig förtrogen med kraven på de olika examensnivåerna.
Tidsbokningsnumret till Vanda tandvård (hammashoito) är (09) 8393 5300.
Du ska teckna en pensionsförsäkring (ArPL-försäkring) (eläkevakuutus (TyEL-vakuutus)) och en olycksfallsförsäkring som omfattar en grupplivförsäkring och en arbetslöshetsförsäkring för de anställda.
Information om studiestödetengelska _ ryska _ estniska _ samiska
Den förälder till barnet som är bosatt i Finland måste vara barnets vårdnadshavare för att barnet ska kunna få uppehållstillstånd.
Du får närmare uppgifter också från tjänsten Studieinfo.fi.
Du kan ta ut högst 18 dagar av din faderskapsledighet samtidigt som barnets mor är moderskaps- eller föräldraledig.
Webbplatsen för sommarteatern Konttisen kesäteatterifinska
Vanligtvis måste du boka en tid hos beskickningen eller tjänstestället i förväg.
Grundnivån är avsedd för personer som kan använda språket i vardagliga sammanhang.
På internet finns en databank för utvecklingsstörda (Kehitysvammahuollon tietopankki) med mycket nyttig information om utvecklingsstörningar och tjänster för handikappade.
Därför får du under dessa dagar inte göra något som kan äventyra ditt tillfrisknande.
Språkcentret vid Lapplands universitet ordnar kurser i finska språket på engelska.
De hjälper dig att integrera dig i Finland.
Du kan få specialvårdspenning från FPA om
Vägledning och stöd för ungafinska _ svenska
Hjälp med fostran av barn
HelMet-biblioteken har en gemensam webbtjänst.
Du kan anlita dessa företag att transportera dina ägodelar från ett land till ett annat och också att packa dina saker och tillhandahålla förpackningsmaterial.
På InfoFinlands sida Tjänster för handikappade hittar du information om tjänster för handikappade.
Jämlikhet på arbetsplatsen
I Finland finns många företag som erbjuder olika typer av Internetanslutningar.
Föreningen har ett resurscenter (voimavarakeskus) i Vanda där man får stöd och råd.
Högre yrkeshögskoleexamina
I Helsingfors och Helsingforsregionen verkar många religiösa samfund.
När du väljer företagsformen ska du beakta bland annat antalet grundare, behovet av kapital, fördelningen av ansvar och beslutsmakt samt finansiering och beskattning.
Vid Stadin ammattiopisto ordnas förberedande utbildning inför yrkesutbildning för invandrare.
Du får mer information om hemkommun på InfoFinlands sida Hemkommun i Finland.
Den gemensamma ansökan ordnas två gånger per år, på våren och på hösten.
Om intyget har utfärdats av en myndighet i ett EU-land och åtföljs av blankett EU 2016/1191, behöver intyget inte översättas.
Kontrollera på förhand vilken typ av avfall stationen tar emot.
Kommunernas finansieringsandelar fastställs utgående från antalet invånare.
Tolkbeställning
när du vill utöka din yrkeskunnighet och dina kunskaper
Du måste dock ha visum eller rätt att vistas i Finland tre månader utan visum.
Mer information om föreningarna hittar du på sidan Vantaalla.info.
Flyktingrådgivningen (Pakolaisneuvonta) ger kostnadsfri juridisk rådgivning till asylsökande, flyktingar och andra utlänningar.
Unga flickor kan söka hjälp vid Flickornas hus som finns på många orter.
Privata jurister och advokater
Om du kommer till Finland för att arbeta behöver du ett uppehållstillstånd.
Hjälp för män att sluta med våldsamt beteendefinska
Information om att köpa en bostadfinska _ svenska _ engelska
När ett barn föds i ett samboförhållande, kan hen få
Du hittar utbildningar på Studieinfo.fi.
I småbarnspedagogiken beaktas familjens religion eller livsåskådning.
Som företagare har du ansvaret för att ge arbetstagarna inskolning i arbetsuppgifterna.
Jourfinska _ svenska _ engelska
Priserna och tjänsterna varierar mycket.
Läs mer om vårdnaden om barn på InfoFinlands sidor Skilsmässa, Familjer med en förälder och Vad är en familj?.
Då utgår man ifrån att båda äger en lika stor andel och denna egendom delas på hälft.
Tolken sköter inga andra uppgifter utöver tolkningen.
Arbetsgivaren har skyldighet att utfärda ett intyg ännu tio år efter att anställningen upphört.
Om du har problem eller oklarheter med uppehållstillståndet, ska du ta kontakt med migrationsverket.
Om du omfattas av den finländska sjukförsäkringen (sairausvakuutus) ersätter FPA (Kela) en del av kostnaderna för många läkemedel.
Adress: Bangårdsvägen 7 (ingång via Loktorget)
Hälsovårdstjänster i Karleby
Kontaktuppgifter till InfoFinlands redaktion:
barnets far är finsk medborgare och föräldrarna är gifta,
Finska är modersmålet för cirka 90 procent av finländarna.
Polisen utfärdar pass för finska medborgare.
Riksdagen utser statsministern och republikens president tillsätter honom eller henne.
Det är viktigt att du ansöker om fortsatt uppehållstillstånd innan ditt tidigare uppehållstillstånd går ut.
När ni överväger att skiljas och behöver hjälp med att komma överens om saker, kan ni ansöka om medling i familjeärenden (perheasioiden sovittelu).
Med papperslösa avses invandrare som inte har uppehållstillstånd eller invandrare som inte har sjukförsäkring.
Om din sjukdom är långvarig och du inte kan arbeta finns det mer information om FPA:s sjukpenning på InfoFinlands sida Stöd när du är sjuk.
NewCo Helsinki ordnar företagarutbildning på finska, engelska och ryska.
Tolken har som uppgift att tolka det som du och myndigheten säger.
Giltigt pass eller annan identitetshandling som styrker ditt medborgarskap
Fortsatt uppehållstillstånd för studerandefinska _ svenska _ engelska
Skyddshemmet Mona är ett skyddshem avsett för invandrarkvinnor och deras barn.
Föreningen har verksamhet i Helsingfors, Tammerfors och Lahtis.
Den unga kan själv ingå ett arbetsavtal.
Försörjningsförutsättningen kan i vissa fall undgås.
Du har rätt att vägra övertidsarbete.
Fråga mer vid din egen hälsostation.
Brådskande reparationer kan dock göras utan ett meddelande.
De största språken efter finska och svenska är ryska, estniska, engelska, somaliska och arabiska.
Om familjens yngsta barn är yngre än tre år kan föräldern få hemvårdsstöd för vård av barnet i hemmet.
Ansök om tillstånd hos kommunens hälsomyndighet innan lokalerna tas i bruk.
I utredningen klarläggs situationen för den sökande och landet där denna kommer ifrån så noga som möjligt.
Om du har problem med att betala räkningar och skulder, kontakta ekonomi- och skuldrådgivningen (talous- ja velkaneuvonta).
Om du har avlagt grundskolan eller gymnasiet utomlands, antas du till en yrkesutbildning enligt prövning.
Genom läroavtalsutbildning kan du avlägga samma examen som vid yrkesläroanstalter.
Om du vill flytta till Finland måste du ha ett uppehållstillstånd eller så måste du
Läs mer på InfoFinlands sida Studerande.
Etableringsanmälan
Du kan ansöka om bidraget vid socialbyrån i din hemkommun.
Vem är asylsökande?
Om du har din hemkommun i Grankulla, kan du utnyttja de offentliga hälso- och sjukvårdstjänsterna.
Du kan söka progressiv beskattning också i efterskott.
På InfoFinlands sida Familjemedlem hittar du mer information avsedd för personer som flyttar av familjeskäl.
På en privat läkarstation måste du betala samtliga kostnader själv.
Kontaktuppgifterfinska _ svenska
På följande villkor:
Läs mer om dessa dagar på sidan Finländska helgdagar.
Du kan be om hjälp i frågor som rör startandet av ett företag hos nyföretagarcentralerna.
Du kan lära dig svenska med hjälp av appar som du kan ladda ned i din telefon eller surfplatta.
Information om dagvården finska _ svenska _ engelska
Du får också ett meddelande när beslutet är klart.
Uppgifternas ämnesområden rör det vardagliga livet såsom fritid, utbildning och vanliga situationer på arbetet.
Huvudregeln är att du omfattas av den sociala tryggheten i Finland och har rätt till FPA:s förmåner om du bor stadigvarande i Finland.
Om du äger en fastighet betalar du vanligen
Du kan söka till många universitetsutbildningar i den gemensamma ansökan till högskolor.
Modern inleder i allmänhet moderskapsledigheten 30 vardagar för det beräknade förlossningsdatumet.
Mer information om upphovsrätt finns på adresserna www.teosto.fi, www.kopiosto.fi, www.gramex.fi, www.tuotos.fi.
Vägledning i högskolestudier
Ofta måste de som arbetar i Finland betala skatt på sin lön till Finland.
Jourmottagningarfinska _ svenska _ engelska
Denna rätt kan inte begränsas med avtal.
Rättshjälp för asylsökande
Länder som är anslutna till Apostilleavtaletengelska _ franska _ spanska _ tyska _ portugisiska
Huvudstadsregionen har goda kollektivtrafikförbindelser.
Inträdesavgifter och rabatter
Om du inte kan återgå till arbetet på grund av sjukdom eller skada kan du ansöka om invaliditetspension (työkyvyttömyyseläke) eller rehabiliteringsstöd (kuntoutustuki).
linkkiRegionförvaltningsverket i Västra och Inre Finland:
Läs mer på InfoFinlands sida Avfallshantering och återvinning.
Äktenskap
Banvägen 2, Dickursby
Barn och unga
Läkaren bedömer situationen.
Dagens stadssund var då en smal havsvik som sträckte sig ända till Kyrkbacken.
Du studerar i gymnasiet
Då minns man de tre vise männen som kom med gåvor till Jesusbarnet.
Läs mer om barnets efternamn på sidan När ett barn föds i Finland.
För omskärelse behövs ett skriftligt samtycke av pojkens vårdnadshavare.
För studerande och förvärvsarbetande lönar det sig att ta reda på om läroanstalten eller arbetsplatsen erbjuder motionsmöjligheter.
Telefon 0295 419 626 tisdag, onsdag och fredag kl. 10.00–11.00
Stadin ammatti- ja aikuisopisto är Finlands största yrkesläroanstalt där man kan utbilda sig inom många olika branscher.
Läs mer på InfoFinlands sida Prövning av hinder mot äktenskap.
I dessa fastställs till exempel minimilöner, arbetstider, semestrar, lön för sjukdomstid och uppsägningsvillkor.
förvärvat kvalifikationer för ett yrke som är reglerat i Finland i ett EU-land, EES-land eller Schweiz,
Kontakta rättshjälpsbyrån om du vill ha ett rättsbiträde.
Intervjuerna görs i de länder där flyktingarna vistas, vanligen i flyktingläger eller i UNHCR:s lokaler.
Stöd och verksamhet för regnbågsfamiljerfinska
din flyktingstatus i Finland har upphört eller återkallats eller det har fattats beslut om att avvisa dig
Mer information hittar du på Esbo stads webbplats.
På biblioteket kan du även låna tidskrifter, e-böcker samt CD- och DVD-skivor.
Information om enskilda jurister finns bland annat på Finlands Advokatförbunds webbplats.
Barnet kan få dispens för att börja i skolan.
Genom att betala en bostadsrättsavgift, som är 15 procent av bostadens anskaffningspris, och därefter varje månad ett rimligt bruksvederlag får man rätt att förvalta över bostaden precis som om den vore en ägarbostad.
Om du är sjuk en lång tid och din arbetsgivare inte längre betalar dig lön under sjukledigheten kan du söka FPA:s sjukdagpenning när lönen inte längre utbetalas.
De måste betala samma avgifter för vården som övriga invånare.
Information om att teckna försäkringar för anställdafinska _ svenska _ engelska
Köpeanbudet är bindande.
Barnets födelseattest om du har vårdnaden om ett barn
Du kan göra brottsanmälan på internet.
Tillfällig hemvård kostar lika mycket för alla.
Du kan meta med metspö och pimpla på isen utan ett separat tillstånd.
Du kan ansöka om underhållsstöd från Fpa i följande situationer:
Du får hjälp på finska och svenska, och på de flesta ställena även på engelska.
När du upptäcker att du är gravid, kontakta mödrarådgivningen eller familjecentret i din hemkommun.
Att börja i skolan
Det är inte obligatoriskt att ange barnets religion.
Migrationsverket beviljar dig fortsatt uppehållstillstånd om grunden för det tidigare uppehållstillståndet fortfarande existerar.
I Finland firas vändagen inte med lika mycket pompa och ståt som till exempel i USA.
Enligt finsk lag är kvinnor och män jämställda.
Etelärinne 32
Om Migrationsverket behöver ytterligare utredningar av dig, meddelas detta i Enter Finland-tjänsten.
Finlands beskickningar utomlandsfinska _ svenska _ engelska
Ryska kejsaren var ändå regent i Finland.
Omskärelse (ympärileikkaus) av flickor är ett brott i Finland. Man kan få ett flera års fängelsestraff för det.
Tvåspråkiga kommuner finns på väst- och sydkusten.
En handikappad har rätt att leva ett vanligt liv, till exempel studera, arbeta och bilda familj.
Bodelning mellan makarfinska _ svenska _ engelska
Hemfrid innebär också att du i regel själv får bestämma vem som har tillträde till ditt hem.
Avlöningsdagen är vanligen en eller två gånger i månaden.
Hyresvärden kräver att jag tecknar en hemförsäkring.
Du behöver eventuellt bifoga till etableringsanmälan också ett utdrag som motsvarar handelsregisterutdraget i Finland, som en myndighet i ditt hemland utfärdar.
Integrationsutbildningen omfattar vanligen studier i finska eller svenska. I utbildningen bekantar du dig med det finländska samhället och arbetslivet och den finländska kulturen.
Trillagatan 5
I Grankulla finns en järnvägsstation och i staden finns många busslinjer.
Icke-medicinsk omskärelse omfattas inte av den offentligt finansierade hälsovården, och kan därför inte göras på en offentlig hälsostation, och man måste själv betala det.
Rehabilitering som ordnas av kommunerna
Du kan inte gå till polikliniken utan en läkarremiss.
är arbetsoförmögen på grund av din sjukdom
Företagsfinland ger upplysningar om olika finansieringsalternativ.
Rådgivning på olika språk:
Högskolor som erbjuder SIMHE-tjänsterfinska _ svenska _ engelska
Läkaren kan vid behov skriva en remiss till ungdomspsykiatriska polikliniken (nuorisopsykiatrian poliklinikka).
Dagvårdsblanketterfinska _ svenska
Män och kvinnor ska behandlas lika vid anställning och beträffande arbetsförhållanden och lönesättning.
Jag har fått för lite lön utbetalad.
Museet för nutidskonst Kiasmafinska _ svenska _ engelska _ ryska
Om du vill byta efternamn ska du meddela detta till magistraten.
Kontaktuppgifter till Marthaförbundetfinska _ engelska
Att ansöka om bostadsbidrag
Invandrare kan även sköta ärenden vid servicestället International House Helsinki.
Uppehållstillstånd för före detta finska medborgarefinska _ svenska _ engelska
Du kan ändå få stöd för den från FPA.
Museer i Helsingforsfinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
När den första ansökan om skilsmässa har lämnats in börjar en sex månader lång betänketid.
Barndagvård
Invandrarenhetenfinska _ svenska _ engelska
Du kan avlägga examen på olika orter i Finland.
linkkiTE-tjänster:
tfn 0400 187 250
Många kliniker har även en jourtid, då man kan komma för vård utan en tidsbokning.
Om du behöver brådskande hjälp av polisen i nödsituationer, ring nödnumret 112.
Information för företagare om företagshälsovårdenfinska _ svenska _ engelska
nivåerna A1 och A2: grundläggande språkkunskaper (peruskielitaito)
Alkoholdrycker är relativt dyra i Finland och köpet av dem begränsas med åldersgränser för unga personer.
På Nuppi kan du till exempel få hjälp med mentala problem och missbruksproblem.
Inträdesprov eller lämplighetsprov ordnas också för många utbildningar.
el och vatten
Äktenskap och uppehållstillstånd
Ta kontakt med en privat läkarstation.
Du kan ansöka om arbets- och folkpension med samma blankett.
Arbetsgivaren ska ordna arbetsplatsintroduktion för nya anställda.
Vilka yrken kan studera till?
Ta med ett intyg över att du omfattas av den finländska sjukförsäkringen.
Den förberedande utbildningen är avsedd för unga och vuxna, som är intresserade av yrkesstudier och vill förbättra sina kunskaper i finska..
Till exempel är tekniska högskolors motsvarighet till magisterexamen diplomingenjörsexamen (diplomi-insinööri).
inkomster
I Finland finns femton ELY-centraler.
svenska 029 497 001
Kom ändå ihåg att arbetsgivaren inte kan ansöka om uppehållstillstånd för dig, utan hen kompletterar din ansökan för egen del i tjänsten Enter Finland.
Jourmottagningen vid Jorv sjukhus
rehabiliteringshandledning
Frivilligarbete är ett bra sätt att hjälpa, lära känna nya människor och medverka i något som du tycker att är viktigt.
Universitetscentret Chydeniusfinska _ svenska _ engelska
Störst är bristen på små bostäder.
Den slutliga beskattningen fastställs utgående från uppgifterna i skattedeklarationen.
Om du inte söker jobb men vill få den inledande kartläggningen och en integrationsplan upprättade, ska du kontakta invandrarenheten vid Helsingfors stads social- och hälsovårdstjänster.
Brottsofferjouren ger även rådgivning för att motarbeta diskriminering.
Det är bra att boka en tid på tjänstestället i förväg.
Till Finland som praktikant
mån–ons kl. 8–16
medborgare i ett nordiskt land och har varit bosatt i Finland de senaste fem åren
Tfn 043 825 0535
På rådgivningen vårdas inte barn som insjuknar plötsligt, men du kan be om råd via den centraliserade telefontjänsten (06) 826 4477.
Tfn (09) 8789 1300
Arbete
Magistraterna lagrar information om invånarna i sitt område i befolkningsregistret.
Som EU-medborgare kan du komma till Finland om du har ett pass eller ett ID-kort förutsatt att du inte har utfärdats ett inreseförbud.
Stöd till arbetslösa invandrarefinska _ svenska _ engelska
Familjemedlem
Kurser i finska språket vid öppna universitetet
Invånarhuset Kivenkolo är ett öppet vardagsum där du kan få rådgivning och handledning på olika språk.
uträtta ärenden,
Hyresbostäderfinska _ engelska
Målet med rehabiliteringen är att hjälpa dig att klara dig bättre i vardagen.
Om du inte företedde en giltig resehandling till myndigheten i samband med din asylansökan får du förvärvsarbeta i Finland när det har gått sex månader sedan du lämnade in din asylansökan.
När du söker till ett vuxengymnasium är inte medeltalet på ditt betyg av betydelse.
Barnpassningsservice för barnfinska _ engelska
Pausen kan vara minst tre månader och högst två år lång.
I gymnasiet läser man samma ämnen som i den grundläggande utbildningen, med undervisningen är mer krävande och studierna mer självständiga.
om utbetalningen av ditt arbetsmarknadsstöd avbryts tillfälligt eftersom du på grund av vården av ditt barn inte kan delta i integrationsåtgärderna eller
Död
Stödets storlek beror bland annat på familjens inkomster och kommunen som familjen bor i.
Fundera noga på om omskärelse behövs.
Du kan även få rabatt på exempelvis olika former av motion och kultur.
Ansökningen kan tas för behandling först när du har besökt beskickningen.
Problem i parförhållandet kan behandlas i par- och familjeterapi.
Ett ofött barns medborgarskap
Du kan anlita vilken som helst rättshjälpsbyrå oberoende av din hemkommun.
Information om den sociala tryggheten för studerandefinska _ svenska _ engelska
Vägledning kan ges individuellt eller i grupp.
tfn 016 322 8091 eller tfn 016 322 8014
Familij
Om du blir arbetslösfinska _ svenska _ engelska
genom ansökan eller anmälan om medborgarskap.
Ett kommanditbolag är ett personbolag som skiljer sig från ett öppet bolag på så sätt att det i kommanditbolaget finns utöver en eller flera ansvariga bolagsmän åtminstone en tyst bolagsman, d.v.s. en person som är delägare i företaget. Vanligen är den tysta bolagsmannen en investerare.
Ange kontonummerfinska _ svenska _ engelska
Den högsta beslutsfattande makten i Karleby stad innehas av stadsfullmäktige.
Socialarbetaren som ansvarar för handikapptjänster i din hemkommun bedömer tillsammans med dig om du behöver göra ändringsarbeten i din bostad.
Socialservicecentret
Också en hemförlossning är möjlig, men den omfattas inte av den allmänna hälsovården och rekommenderas inte.
FPA-kort
Det är bra att anlita en jurist för upprättandet av bouppteckningen.
Behöver du en jurist?
I Karleby finns grupper för den förberedande utbildningen i lågstadiet i Hollihaan koulu och Koivuhaan koulu och i högstadiet i Stenängens skola.
Du kan också ha rätt till den sociala tryggheten i Finland om du arbetar i Finland.
Tjänsten är avsedd för personer som har bristfälliga kunskaper i finska, svenska eller engelska.
linkkiHelsingfors kyrkliga samfällighet:
ditt uppehållstillstånd inte begränsar vilken arbetsgivare du får arbeta för
Fpa betjänar sina kunder på sina byråer, per telefon och post samt via webbtjänsten som finns på FPA:s internetsidor.
Med hjälp av dem kan du på förhand uppskatta om du kan betala tillbaka lånet.
Esbo stad ordnar mycket verksamhet för de föräldrar som vårdar barn i hemmet. Det finns till exempel invånarparker, öppna daghem och klubbar.
Rätt att få eget sjukförsäkringskort.
Information till en avlidnes anhörigfinska _ svenska
Mer information om resekorten och deras försäljningsställen i Esbo hittar du på HRT:s webbplats.
Aktiveringsmodellen för arbetslöshetsförsäkringen finska _ svenska _ engelska
Betalningen av dagpenning inleds efter en självrisktid (omavastuuaika).
Källskattekort måste du ansöka med en pappersblankett.
Du får vistas i Finland eller något annat land i Schengenområdet utan uppehållstillstånd så länge som ditt visum är i kraft.
Thai
De flesta invånarna i Rovaniemi äger sin bostad. De har tagit lån eller finansierat sin bostad på andra sätt.
Om du har bokat en tid hos tandläkaren, men inte kan komma på avtalad tid ska du komma ihåg att avboka din tid.
intyg på studier i tjänstemannafinska eller -svenska som du har avlagt vid universitet eller högskola
På cykel och till fots
Medicinsk rehabilitering kan ordnas i ett rehabiliteringscenter eller som öppen terapi. Under den öppna terapin kan du bo hemma.
Barn med invandrarbakgrund och barn från tvåspråkiga familjer kan få hemspråksundervisning (oman äidinkielen opetus) om tillräckligt många barn anmäler sig till gruppen för det egna språket.
Prövotiden kan vara högst sex månader.
Betala samtidigt också ansökningens handläggningsavgift.
Parktanterna erbjuder tillfällig hjälp med skötsel av barn på förmiddagar.
Seniorernas hälsopunkterfinska _ svenska
Ett öppet bolag bildas då två eller fler personer kommer överens om att grunda ett bolag genom att teckna ett bolagsavtal.
Simhallar
Registrerat parförhållande
Anslutningarnas priser varierar mycket.
Arbetsmarknadsstödet är behovsprövat, vilket betyder att dina andra inkomster och din situation som en helhet påverkar dess belopp.
linkkiCentralen för främjande av Folkmusik och Folkdans :
På turistbyrån finns bland annat broschyrer om Rovaniemi, kartor, tidtabeller och information om evenemang.
Ibland kan det utöver dessa förekomma övriga villkor.
En arbetstagare är skyldig att
Ofta behövs ett domstolsbeslut för utmätning.
Det firas på självständighetsdagen den 6 december.
Information om olika sätt att delta och påverka finns på stadens webbplats.
Då hanteras plötsliga sjukdomar och olyckor vid jouren.
Hyra betalas vanligen en gång per månad.
Om du vill hyra en privat hyresbostad ska du kontakta den som hyr ut bostaden. Kom överens om när du kan gå och titta på bostaden.
Att ansöka om finskt passfinska _ svenska _ engelska
Hjälp för män
Ansökan om uppehållstillstånd är avgiftsbelagd.
På MoniNets webbplats finns en studiemiljö för finska språket där du kan studera finska på egen hand.
Med freden etablerades den katolska tron i Finlands västra delar och den ortodoxa tron i landets östra delar.
Juridisk rådgivning till brottsofferfinska _ svenska _ engelska
Fråga din arbetsgivare som hen använder tjänsten Enter Finland för arbetsgivare.
Adoption inom familjen betyder att makan/maken adopterar sin makas/makes barn och blir officiellt barnets andra förälder.
du omfattas av den sociala tryggheten i Finland.
Folkhögskolorna ordnar vanligen två olika slags undervisning, kortkurser (lyhytkurssi) och långa utbildningslinjer (pitkä opintolinja).
Om du är orolig för en närstående person och tror att han eller hon kan vara i behov av hjälp, kan du rådfråga till exempel hälsovårdaren eller läkaren vid hälsocentralen.
Om tiden inte passar ska du ringa tidsbokningen och boka om tiden.
Tfn (09) 4716 7060
Finsk konst presenteras till exempel i Ateneum som hör till Nationalgalleriet och Esbo moderna konstmuseum (EMMA). Med
Kommunernas rehabilitering omfattar:
Tolknings- och översättningstjänsterfinska _ svenska _ engelska
När ska jag betala hyresdepositionen?
Där hittar du även kontaktuppgifterna till beskickningarna.
Läs mer på InfoFinlands sida Ekonomiska problem.
Tfn (09) 81621
familjens inkomster
SERI-stödcentretfinska _ svenska _ engelska
VAR: röda batteriinsamlingslådor i butiker och kiosker
Tandvården vid hälsovårdscentralen är kostnadsfri för barn under 18 år.
Utkomstskydd för arbetslösa
Du får:
barnfamiljer
På språkkaféerna samtalar man på finska, så det är bra om du redan kan lite finska.
Hos en privat tandläkare måste du betala samtliga kostnader själv.
I staden finns även möjlighet till mångkulturell dagvård, familjedagvård och specialdagvård.
ta torra eller kullfallna träd, ris, mossa eller liknande på annans mark utan tillstånd
Bodelningsmannen tar betalt för arbetet.
Om du vill ha kontakt med en anhörig som försvunnit kan du be om hjälp vid personefterforskningen vid Finlands Röda Kors.
Karleby stad grundade museet 1909 utgående från en testamentsgåva av affärsmannen Karl Herman Renlund (1850–1908) .
För den som säljer en fastighet varar ansvaret fem år.
I stora städer kan könssjukdomar vårdas på polikliniker för könssjukdomar (sukupuolitautien poliklinikka).
På webbplatsen för föreningen för familjer med en förälder, Yhden Vanhemman Perheiden Liitto ry, finns information och råd för föräldrar som överväger skilsmässa.
däck
Om tandvården för barn under skolåldern får du information på barnrådgivningen (lastenneuvola) och vid tandklinikerna (hammashoitola).
När du fyllt i anmälan, kom ihåg att följa ditt konto i tjänsten Enter Finland.
Mer information finns på tjänsten HelsingforsRegionen.fi.
Du ansöker om lånet i banken när du har fått FPA:s beslut om statsgaranti.
Kollektivtrafikfinska _ svenska
Skriv ut blanketten på Migrationsverkets webbplats och fyll i den färdigt.
Efter utgången av moderskapspenningperioden kan en av vårdnadshavarna ta ut föräldraledighet.
På de största orterna finns flera privatläkare och på somliga orter också privata rådgivningsbyråer.
Om du har flera arbetsgivare
Att grunda en förening
I Helsingfors finns många bibliotek på olika håll i staden.
NewCo Helsinki ordnar företagarutbildningar på finska, engelska och ryska.
Från studerande till anställd
Om du studerar vid gymnasium, yrkesläroanstalt, yrkeshögskola eller universitet kan du söka bostad hos Domus Arctica-stiftelsen.
Också dina familjemedlemmar kan ha rätt till dessa tjänster om de flyttar till Finland tillsammans med dig.
Tandläkarjouren (kvälls-, vardags- och helgjour) ordnas vid polikliniken för tand- och munsjukdomar vid Mellersta Österbottens social- och hälsovårdssamkommun Soite, Mariegatan 16–20, 67200 Karleby (vån 1, del D), vardagkvällar kl. 16.00–21.00 samt veckoslut och helgdagar kl. 8.00–21.00.
En ung i åldern 13–22 år kan få hjälp vid Ungdomspolikliniken Nupoli om hen har problem till exempel med den mentala hälsan, rusmedelsbruk, spelande eller fritidsaktiviteterna.
Bibliotek
Undervisningstillståndfinska _ svenska
Där hjälper experterna dig att utveckla affärsidén, göra en marknadsundersökning, beräkna lönsamheten och kartlägga finansieringen.
Då bostadsbidraget kalkyleras avsätts 300 euro per månad av dina förvärvsinkomster.
Du kan be bibliotekarien på ditt eget bibliotek att beställa det material du vill ha åt dig.
Till exempel inom social- och hälsovårdsbranschen fattas beslutet av Valvira, och inom undervisningssektorn av Utbildningsstyrelsen.
Det är viktigt att kunna diskutera konflikterna inom familjen.
Du kan också behålla ditt eget efternamn eller ta ett dubbelnamn.
I ett samboförhållande kan makarna ha ett gemensamt efternamn.
Om tjänsten är hårt belastad, kan du lämna ett meddelande om att bli uppringd vid ett senare tillfälle.
Ett tidsbestämt hyresavtal får inte sägas upp under dess löptid.
Startpunkten i Iso Omena
Magisterprogrammen pågår i cirka två år.
Du kan också söka dagvårdsplats via Internet.
När du letar efter en bostad är det bra att räkna med att det tar till och med flera månader.
Läs mer: Graviditet och förlossning.
Hälsovägen 4
Magistraten i Lappland
Information om VALMA-utbildningarfinska
Rovala-institutets utbildning för invandrare
Information om social trygghetfinska _ svenska _ engelska
Skatteåterbäringen betalas antingen direkt på ditt bankkonto.
Läs mer linkkiFörsamlingen:
Bastu, tvättstuga och bilplats
Då är den unga en myndig samhällsmedlem som har rätt att besluta om sitt eget liv.
Läs mer: Att grunda ett företag
främjande av invandrares integration
Kunta-asunnot Oy:s bostäder
Finland är en av de bästa länderna i världen om man vill se norrsken (aurora borealis).
Utbildningen kan vara till exempel studier i finska eller yrkesutbildning.
Att ta sig till arbetet eller butiken till fots eller med cykeln är ett lätt sätt att få den dagliga motionsdosen.
De vuxna i familjen kan vara av samma eller olika kön.
Grunden för diskriminering kan vara till exempel etniskt ursprung, nationalitet eller religion.
uppdrag inom företagsledning
Ruttjänstenfinska _ svenska _ engelska
Ansvaret för skötseln av barnen och hemmet hör till både kvinnan och mannen.
de skatter som har betalats på dina inkomster från början av året
Du kan teckna en försäkring hos ett försäkringsbolag i ditt hemland eller fråga om en lämplig försäkring hos internationella försäkringsbolag.
Mer information om sådana situationer får du vid FPA.
På vissa orter utkommer även svenskspråkiga tidningar.
Dina möjligheter att få en bostad påverkas av ditt bostadsbehov och dina tillgångar och inkomster.
Ansök om moderskapsunderstöd och moderskapspenning hos FPA senast två månader före det beräknade förlossningsdatumet.
Finlands röda kors (FRK) hjälper kvotflyktingar när de flyttar till Finland.
I Karleby finns nära på hundra idrottsföreningar för olika grenar samt föreningar som arrangerar övrig motion.
Övriga studiemöjligheter
Sexuellt våld kan även förekomma i parförhållanden och äktenskap.
samma uppgifter för de personer som har rätt att använda kontot.
Flygplatsenfinska _ svenska _ engelska _ ryska _ kinesiska
Om du blir sjuk eller skadas, har du rätt till brådskande vård inom den offentliga hälso- och sjukvården, till exempel på en hälsostation eller ett sjukhus.
Med grundlagen stadgas till exempel de grundläggande rättigheterna för alla som är bosatta i Finland samt regler för hur den finska staten fungerar.
Sammanlagt väljer man 200 riksdagsledamöter.
Vid vuxengymnasiet är studierna flexibla.
Du hittar kontaktinformation på Global Clinic:s hemsidor.
Tfn 09 276 62 8 99
Om du har hemkommun i Finland får du sjukvården förmånligare.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
I våldssituationer får du mer information på InfoFinlands sida Våld.
Om föräldrarna inte är gifta, får barnet finskt medborgarskap av sin far enligt följande:
arbetsplats eller eget företag i Finland
Tfn 029 5660 160
Det är också bra att nia äldre människor.
Alla har rätt till företagshälsovård
i något annat religiöst samfund som är registrerat i Finland.
Information om grannmedlingfinska _ engelska
Allmän information om studier i finska och svenska i Finland hittar du på InfoFinlands sida Finska och svenska språket.
Även samkönade par kan gifta sig i Finland.
På detta inverkar om du flyttar till Finland från
Du kan till exempel ersättas med en felfri vara eller få dina pengar tillbaka.
I den privata sektorn kan arbetsgivaren själv bedöma huruvida den anställdas utländska examen godtas.
Rådgivningstjänsterna i den egna hemkommunen är gratis.
Du kan söka sjukdagpenning om du:
Boende
När du köper en bostad måste du också betala överlåtelseskatt (varainsiirtovero).
adress i Finland eller i ett annat land
De har ofta öppet också på kvällarna och ibland får man fortare en tid där.
Alexandersgatan 9 (Gloet)
Tolkningen kan också ordnas per telefon.
Hela saker är inte avfall.
Om ditt äktenskap eller registrerade parförhållande upphör
Om barnets sjukdom inte kräver omedelbar vård ska du vänta tills din hälsostation har öppet igen.
Om du vill avlägga en fristående examen ska du ta kontakt direkt med läroanstalten.
Byggherrarnas kontaktuppgifterfinska
Kommunen ska dock säkerställa att invånaren har råd med att bo i ett servicehus om han eller hon är i behov av serviceboende.
Väg in i arbetslivet
En jurist svarar på dina frågor till exempel om arbetsavtal, lön eller arbetstider.
Förbered dig på företagande genom att skaffa så goda kunskaper och färdigheter som möjligt, eftersom det är riskabelt att starta ett företag utan tillräckligt kunnande och tillräckliga språkkunskaper.
Information om begravning får du på Vanda församlingars gravkontor (Vantaan seurakuntien hautaustoimisto) och vid privata begravningsbyråer (hautaustoimisto).
dagtid kl. 8–22
Kurserna är avgiftsbelagda.
I Esbo finns även Vi läser tillsammans-grupper, där kvinnor kan studera finska språket.
Du kan ansöka om permanent uppehållstillstånd på internet i tjänsten Enter Finland.
Förskoleundervisning ges på finska och på svenska.
Om du har bett om ett arbetsintyg men inte fått det, ska du kontakta arbetarskyddsmyndigheterna.
Tfn (09) 83 911.
Stenbäcksgatan 9
Den är öppen mån-tors kl. 8–15 och fre kl. 8–13.
Sveriges kung Gustav Vasa grundade Helsingfors på stranden av nuvarande Gammelstadsforsen genom att den 12 juni 1550 beordra invånare i andra städer att flytta till Helsingfors.
Mer information om barnskyddet finns på InfoFinlands sida Barnskydd.
I kallelsen anges tolkningsspråket, den exakta adressen till verksamhetsstället där samtalet hålls och klockslaget.
Förbund för studerande vid yrkeshögskolorfinska _ svenska
Den som bor i en stödbostad klarar nästan självständigt av de dagliga bestyren.
Om du är sjuk en lång tid och din arbetsgivare inte längre betalar dig lön under sjukledigheten kan du söka FPA:s sjukdagpenning när lönen inte längre utbetalas.
Ordbok i det finska teckenspråketfinska
Är ett muntligt avtal tillräckligt?
Länkar till kommunsidorna hittar du med hjälp av Menyn Städer i höger spalt.
tfn 016 328 2100
Mer information hittar du på Nödcentralsverkets webbplats.
Peliklinikka
För progressiv beskattning behöver du ett skattekort för begränsat skattskyldiga (rajoitetusti verovelvollisen verokortti).
Information om den inkomstrelaterade dagpenningenfinska _ svenska _ engelska
Servicepunkter finns på olika håll i staden.
När ett barn insjuknar - råd till föräldrarnafinska _ svenska _ engelska
kollektivavtalet som tillämpas på arbetet
I Rovaniemi stad finns 23 skolor med årskurserna 1–6, Lapplands övningsskola som upprätthålls av
Vid kallt väder lönar det sig att ha på sig flera lager med kläder.
Du kan också kontakta en läroanstalt som tillhandahåller läroavtalsutbildning.
Ansökan ska lämnas in senast inom tre månader från datumet för inresa.
Vid högskolornas SIMHE-tjänster kan du söka hjälp och information om högskoleutbildning i Finland och om hur du ansöker till högskoleutbildning.
Mervärdesskattebeloppet varierar emellertid för olika produkter.
Också före detta finska medborgare räknas som återflyttare.
Mer information får du på InfoFinlands sida Företagshälsovården och på social- och hälsovårdsministeriets webbplats.
Det finns ofta en bastu i finländska hem.
Mer information om ämnet hushåll finns på InfoFinlands sida boende.
Kommunen övervakar också den privata dagvården.
Detta betyder att sexuellt umgänge med barn under 16 år är straffbart. (Undantag från detta är en sexuell förbindelse mellan två ungdomar som befinner sig på samma utvecklingsstadium.)
evangelisk-lutherska kyrkan (evankelis-luterilainen kirkko)
Nämnden behandlar inte diskrimineringsfall förknippade med arbetsförhållanden.
Efter tre års boende tryggar dock garantipensionen ett existensminimum.
Hos företagsrådgivningen kan du få hjälp med frågor kring företagets verksamhet eller utveckling.
Arbets- och näringsbyrån stöttar dig i jobbsökningen
Med ett identitetskort för utlänningar kan du styrka din identitet i Finland.
Kristi himmelsfärdsdag
I InfoFinland hittar användaren pålitlig information på sitt eget språk om flytten till Finland, arbete, studier, boende, utbildning, hälsa, familj, problematiska situationer och fritid.
Rådgivningsbyråernas kontaktuppgifterfinska _ svenska _ engelska
Skolveckan består av ungefär 20 lektioner.
Tfn (09) 310 5018 / 116 117
Arbete under moderskapsledigheten är tillåtet om det kan utföras utan att moderns, fostrets eller barnets säkerhet äventyras.
du har fyllt 20 år
På de flesta arbetsplatser är det nödvändigt att kunna finska.
Jämlikhet och jämställdhet i arbetslivet
För att få FPA:s bidrag för psykoterapi ska terapeuten ha rätt att använda psykoterapeutens yrkesbenämning och vara godkänd av FPA.
Tfn 09 839 32622, 09 839 27525 eller 09 839 31766
Det finns skäl att förbereda dig omsorgsfullt för inträdesprovet.
Ett registrerat parförhållande upplöses på samma sätt som ett äktenskap.
ett deltidsarbete, i genomsnitt högst 25 timmar per vecka under terminen
Läs mer: Flytta till Finland.
På InfoFinlands sida Ansökan till utbildning hittar du information om hur du ansöker som examensstuderande till gymnasier, yrkesläroanstalter eller högskolor i Finland.
Den förberedande utbildningen är avsedd för unga och vuxna som vill studera vid gymnasium men saknar tillräckliga språkkunskaper för gymnasiestudier.
Invandrare och grundskolan
Den underhållsskyldiga föräldern har inte betalat det bekräftade underhållsbidraget (Fpa indriver det hos denne senare).
Han eller hon har också rätt att träffa den förälder som han eller hon inte bor med.
Innehållet i yrkesinriktad arbetskraftsutbildning varierar mycket.
Du kan ta dig till ett skyddshem om det på grund av våld är för farligt att vistas hemma.
Småbarnspedagogik.
Förgiftningar, vård och förebyggande: (09) 471 977
Läs mer: Sexuell hälsa.
Du kan besöka Global Clinic även om du inte behöver brådskande sjukvård.
På InfoFinlands sida Missbruksproblem hittar du information om var du kan få hjälp om du eller en närstående till dig har problem med rusmedel.
Boka en tid vid tjänstestället.
Läs på InfoFinlands sida Arbets- och näringsbyråns tjänster vad som krävs för att du ska kunna bli kund hos arbets- och näringsbyrån.
När ett barn föds till familjen har föräldrarna rätt att ta familjeledighet, det vill säga stanna hemma för att ta hand om barnet.
Om du har omskurits innan du kom till Finland och planerar graviditet, kan du låta operera dig för att få slidmynningen öppnad (avausleikkaus).
Båda föräldrarna kan inte vara föräldralediga samtidigt.
Negativt beslut
Båda makarna ska underteckna äktenskapsförordet och två vittnen ska vidimera underskrifterna.
Uppehållstillstånd (om du behöver uppehållstillstånd i Finland)
Man kan ansöka om en plats inom den kommunala dagvården året runt.
Man kan även lämna in bostadsansökan på papper.
Regionförvaltningsverkenfinska _ svenska _ engelska
_ holländska _ rumänska _ ungerska _ italienska
I allmänhet får du nycklarna till bostaden när du betalat hyresgarantin.
Kontaktuppgifter till den landsomfattande telefontjänsten finska _ svenska _ engelska
Giftinformationscentralens telefontjänst är öppen 24 timmar om dygnet. Telefonnumret är (09) 471 977.
Bostadslöshet
Hjälp till brottsofferfinska _ svenska _ engelska
Arbetsgivaren kan lämna uppgifterna om arbetet och sitt företag själv samt följa handläggning av ansökan direkt via tjänsten Enter Finland.
linkkiMedborgararenan:
Permanent uppehållstillståndfinska _ svenska _ engelska
Lagstiftning som rör barn, unga och familjerfinska _ svenska _ engelska
Stadens ungdomsgårdar är öppna för alla ungdomar i åldrarna 10–17 år.
Om du tar med dig en bil till Finland måste du registrera den och betala bilskatt (autovero) för den innan du kan använda den i trafiken.
mån kl. 9–16 utan tidsbeställning
Fortsatt uppehållstillstånd
Barnet får specialundervisning om det har inlärnings- eller koncentrationssvårigheter.
Biblioteket är en plats där du kan låna böcker, läsa tidningar, använda datorn, studera eller delta i olika evenemang.
PB 1
Dessa människor arbetar till exempel i följande arbetsuppgifter:
Tjänsten ger även råd om beskattningen för personer som kommer från utlandet till Finland för att arbeta och skyldigheterna för dem som betalar skatter i internationella sammanhang.
Elektronisk tidsbeställningfinska _ svenska _ engelska
Om du behöver brådskande hjälp av polisen i en nödsituation, ring nödnumret 112.
Du kan också köpa ett prepaid-abonnemang.
Barnbidrag betalas ut månatligen antingen till moderns, faderns eller en annan vårdnadshavares bankkonto.
I verksamheten ingår lek och ledda aktiviteter, till exempel musik, motion och utflykter.
Verksamhet och evenemang för ungafinska _ svenska _ engelska
Väestöliitto ger råd till invandrarfamiljer i frågor rörande barnfostran och familjens välmående.
Om du flyttar till Finland för att bo här stadigvarande i ett år eller längre, ska du också registrera dig i magistraten på din hemort.
Vissa myndigheter godkänner även handlingar på andra europeiska språk.
Under dessa dagar kan modern inte vara moderskapsledig samtidigt.
Om du behöver hjälp och stöd för din mentala hälsa kan du boka en läkartid vid hälsostationen.
Om du är en före detta finsk medborgare kan du återfå ditt finska medborgarskap genom att göra en medborgarskapsanmälan (kansalaisuusilmoitus).
Ring inte nödnumret om det inte är en brådskande nödsituation.
Mer information om myndigheterna och deras uppgifter hittar du på InfoFinlands sida Viktiga myndigheter.
Du kan högst ta ut ett visst maximibelopp.
Lapplands landskapsmuseumfinska
Om du upplever att du behandlats fel inom hälsovårdstjänsterna ska du först reda ut situationen vid din egen vårdenhet.
Hur stora vårdkostnader som försäkringen måste täcka beror på hur länge dina studier varar.
Du kan studera mindre än 90 dagar i Finland utan uppehållstillstånd.
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
Om du inte är säker på om du har hemkommun i Finland kan du ta reda på din situation vid magistraten (maistraatti).
Ansökan till yrkesutbildning i den gemensamma ansökanfinska _ svenska
Bibliotekskortet är avgiftsfritt.
Tfn (09) 4711
Vid behov hjälper mottagningscentret dig.
linkkiFreelanceri.info:
Vaccinationerna är frivilliga.
Det är bra att anlita en kunnig jurist för upprättandet av avtalet.
Startpengen beviljas av den TE-byrå där du är kund.
Alla har rätt till likabehandling.
Krismottagningfinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Kontakta arbetsgivarna direkt
Tfn (09) 276 62899
Man ansöker om skilsmässa med en skriftlig ansökan.
Läs mer: Arbetslöshetsförsäkring.
Tjänsterna hos privatläkare är mycket dyrare för klienten.
Uppsägningstiden för hyresgäster är en kalendermånad.
Skatteprocenten räknas på inkomsterna för hela året.
Att skaka hand är ett vanligt sätt att hälsa på människor i officiella situationer.
Äktenskapsförordet är frivilligt.
I nödfall, om du till exempel inte har pengar för mat, kan du även kontakta diakoniarbetaren i din församling.
I Finland finns ett frivilligt system med arbetslöshetskassor.
Ombudsmannen kan även vid behov be den som misstänks för diskriminering om en redogörelse för det skedda.
Äktenskap mellan två personer av samma kön har varit tillåtet i Finland sedan 1.3.2017.
Om du blir antagen till yrkeshögskolan behöver du inte avlägga de kurser som du redan har avlagt vid öppna yrkeshögskolan.
Om du vill att ditt barn ska få en vaccination som inte ingår i vaccinationsprogrammet ska du beställa tid till en läkare.
Lediga jobb
Utländsk examen i Finland
Ofta ska du själv ingå ett elavtal.
Du kan söka privata hyresbostäder i Esbo via hyresvärdarnas webbplatser:
Bästa stället att fråga mer om kommunernas idrottsplatser är vid idrottsväsendet i den egna kommunen.
I detta fall betjänas du ofta av ditt hemlands beskickning i något av Finlands grannländer.
Barn, vars modersmål inte är finska eller svenska, studerar finska eller svenska som andraspråk i den så kallade S2-undervisningen.
Överlåtelseskatt
Hemförsäkringen kan eventuellt ersätta hyran för en tillfällig bostad.
Information om skolhälsovårdenfinska _ svenska _ engelska
Många vuxengymnasier erbjuder finskakurser för invandrare.
En förening bör inte grundas i syfte att idka en näring.
Du kan använda tjänsterna vid rådgivningsbyrån eller familjecentret om du har en hemkommun i Finland.
I vissa branscher finns också andra obligatoriska försäkringar.
I Furumo i Vanda finns dessutom Vandas och Helsingfors gemensamma begravningsplats för avlidna personer som inte har varit medlemmar i något religionssamfund.
Några gånger per år lottar vi ut priser bland alla som svarat.
Du får skattenumret från skattebyrån samtidigt som du går efter skattekortet.
Arbetsgivaren ska utarbeta ett verksamhetsprogram för arbetarskyddet (työsuojelun toimintaohjelma) som tar upp de säkerhets- och hälsorelaterade riskerna på arbetsplatsen och hur man undgår dem.
För en utvecklingsstörd person finns olika slags specialtjänster.
Hyresbostäder enligt stadsdelfinska _ svenska
Vid folkhögskolan kan du utbilda dig till ett yrke.
Du har tillstånd att:
Den unga kan ställas till svars för brott som han eller hon begått.
Om föräldrarna har olika efternamn beror barnets efternamn på situationen.
Registrering av föreningen
Alla som bor eller vistas i Finland måste följa Finlands lag.
En borgerlig vigsel är avgiftsfri om den sker i magistratens eller tingsrättens lokaler under tjänstetid.
I Esbo finns ungdomsgårdar med utbildade ledare som övervakar verksamheten.
gymnasiet studentexamen
Mentalvårdstjänsterfinska _ svenska _ engelska _ ryska
hemvårdare eller barnskötare.
Väestöliittos karriärmentorskap är avsett för utbildade invandrare.
Information om våld i familjen eller parförhållandet hittar du på InfoFinlands sida Våld.
på finska: 0295 020 701
Seniorrådgivningen
Innehållet i yrkesinriktad arbetskraftsutbildning varierar mycket.
Evenemang och platser i Helsingforsfinska
tfn 016 328 2140
Privata hälsovårdstjänsterfinska
När du flyttar till Finland ska du besöka magistraten (maistraatti)på orten där du är bosatt.
Festivaler i Finlandfinska _ svenska _ engelska _ ryska _ franska _ kinesiska _ tyska _ japanska
Läs mer om språkstudier i InfoFinlands avsnitt Finska och svenska språket.
Hyresvärdens uppsägningstid beror på hur länge hyresavtalet varit i kraft.
Han eller hon tolkar det som du och myndigheten säger.
Studentskrivningarna ordnas på våren och på hösten.
Att ansöka om en bostadsrättsbostadfinska _ svenska _ engelska
När du ansöker om medborgarskap, bifoga ett intyg över dina språkkunskaper.
EU-medborgare som har sin hemkommun i Finland kan rösta i val till Europaparlamentet i Finland om de har anmält sig till rösträttsregistret.
Även då måste hen försöka i förväg komma överens om detta med dig.
på svenska och engelska tfn +358 (0)20 692 226
Det är bra att klarlägga med arbetsgivaren vilka försäkringar han eller hon har tecknat åt sina anställda.
Det kan vara bra att lära sig finska eller svenska trots att du inte tänker bo en lång tid i landet.
Tolktjänster för handikappadefinska _ svenska
Utbildning skattas högt i Finland och det är viktigt att föräldrarna uppmuntrar skolgången.
Eleverna kan själva besöka hälsovårdarens mottagning om de har problem.
ha kvar era egna efternamn eller
Information om körkortfinska _ svenska
Du har rätt att arbeta tills du har fått ett lagakraftvunnet beslut på din asylansökan.
Inomhusmotionfinska _ svenska _ engelska
Då är tolkningen avgiftsfri för dig.
Tfn 020 634 0200 (finska och engelska), 020 634 0300 (svenska)
Man ansöker till förskoleundervisningen med en elektronisk blankett.
Om en av dina familjemedlemmar, som flyttar med dig till Finland, inte är medborgare i ett nordiskt land, kan han/hon behöva uppehållstillstånd eller ett registreringsintyg över uppehållsrätt för EU-medborgare.
skogsvårdsarbete
Boka tid för vigseln hos magistraten.
Den förberedande undervisningen är avsedd för 6-åriga barn med invandrarbakgrund.
TE-byråns tjänster
Du ansöker om hemvårdsstödet hos FPA.
Tfn (09) 310 49999.
När barnet är fött kan faderskapet fastställas hos barntillsynsmannen i hemkommunen.
Om du har ett handikapp eller en sjukdom som försämrar din funktionsförmåga sammanhängande under minst ett år kan du få handikappbidrag (vammaistuki).
Familjehusfinska _ svenska _ engelska
Om du inte gör rättelserna i webbtjänsten MinSkatt, hämta pappersblanketter för rättelserna på Skatteförvaltningens webbplats eller i skattebyrån.
företagsinkomst
Du ska anmäla dig till kursen i förväg: fyll i anmälningsblanketten, lämna den till Rovalas kontor och betala kursavgiften.
Naturen är som bäst en källa till kraft och inspiration.
Fakta om diabetesfinska _ svenska
Om du arbetar i Finland längre än tre månader måste du ansöka om uppehållstillstånd.
Till Finland på grund av familjebandfinska _ svenska _ engelska
att man söker sig till en utbildning på basis av sin utländska utbildning
Du kan själv bestämma om du tar ut hela faderskapsledigheten eller bara en del av dagarna.
Färdtjänst och följeslagartjänstfinska _ svenska
Grundskolan är gratis.
Broschyren Barnets rättigheterfinska _ svenska _ engelska _ ryska
Vid alla hus finns inte alltid samtliga insamlingskärl.
Övriga länder
Först lämnar man in skilsmässoansökan.
Att ansöka om yrkesinriktad rehabiliteringfinska _ svenska _ engelska
Du kan ansöka om uppehållstillstånd för företagare eller uppehållstillstånd för uppstartsföretagare på internet via tjänsten Enter Finland.
Privat tandvård är dyrare än offentlig tandvård.
Du kan ordna säkerheten till exempel så att
Till exempel beaktas inte royaltyn och anställningsoptioner vid beräkning av dagpenningens belopp.
Information för könsminoriteterfinska
Om du behöver en tolk för den inledande kartläggningen och integrationsplanen, måste myndigheten beställa en tolk.
Webbappen IHH Service Advisor App hjälper dig att hitta rätt myndigheter och i den hittar du information om vilka dokument du ska ta med på besöket.
på svenska, tfn 029 502 4881
Information om Finlandengelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
Hyresvärden kan säga upp hyresavtalet om du inte klarar tillräckligt många kurser.
Ungdomsarbete
Det slutliga bostadsbidraget beräknas på följande sätt:
Familjerådgivningens tjänster är konfidentiella och avgiftsfria.
Finskan har färre prepositioner än till exempel de indoeuropeiska språken.
Ohjaamos personal hjälper dig om du inte har ett arbete eller en studieplats.
Lämna blanketten till den lekpark som anmälan i första hand gäller.
Största delen av dessa utbildningar är avsedda för vuxna.
I kommunen finns en socialarbetare som ansvarar för tjänsterna för handikappade.
linkkiAteneum:
Du kan även be om råd gällande andra saker, till exempel boende och ekonomi.
Familjerådgivningarfinska _ svenska
Mun- och tandhälsovårdenfinska _ svenska
Om du är studerande kan du få en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS.
köra ett motorfordon i terrängen utan tillstånd av markägaren
Vaccinationerna ges på barnrådgivningen (lastenneuvola) och inom skolhälsovården.
Utländska studerande får vanligen inget studiestöd.
Specialvårdspenning
säga upp och häva ett arbetsavtal inom ramen för begränsningarna i lag
I juridiska ärenden får du hjälp av en jurist.
Information om hemspråksundervisningfinska
Lapplands yrkesinstitut
Blanketten får du på utrikesministeriets webbplats och från beskickningar i Schengenländer.
I Vanda finns sju hälsostationer (terveysasema) som tillhandahåller offentliga hälsovårdstjänster.
Avfallshantering och återvinning
Moderskapsledigheten är 105 vardagar.
TE-byrån undersöker uppgifterna som du lämnar.
Du behöver inte betala för tjänsterna vid rådgivningsbyrån.
Ungdomstjänsterfinska _ svenska _ engelska
Yrkeshögskolor
Utbildning för invandrare
När du behärskar språket är det lättare för dig att trivas i landet och anpassa dig till livet i Finland.
Våld
Läs mer: Missbruksproblem.
Brandsäkerhet
Flyktinghjälpen hjälper flyktingar och invandrare till exempel i frågor som rör integrationen, boendet och grundandet av egna organisationer.
Stadens hyresbostäder förvaltas av Espoon Asunnot Oy (Espoon Asunnot Oy).
I Vanda finns flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
Också flyktingens familjemedlemmar kan få uppehållstillstånd i Finland.
Om du behöver akut tandvård på en vardag, ska du ringa tidsbokningen så fort den öppnar.
Simhallen i Korso har ett eget simpass för invandrarkvinnor och -flickor.
Erkännande av yrkeskvalifikationer som förvärvats i ett EU-landfinska _ svenska _ engelska
linkkiFinlands Begravningbyråers Förbund:
Vanligtvis måste du boka en tid hos beskickningen i förväg.
Människor som återhämtar sig från problem med den mentala hälsan och missbrukarproblem
Också kännedom om de egna kunderna och försäljningsmetoderna är viktig.
Arbetsgivaren får inte fråga om din familj, vilken religion du har eller om du är politiskt aktiv.
Innan dess kunde två personer av samma kön endast ingå ett registrerat partnerskap.
Serviceställets kontaktuppgifter:
Det är även diskriminering att skapa en hotfull, fientlig, nedsättande eller förödmjukande atmosfär.
Om din bostad har skadats
Kontaktuppgifterfinska _ svenska _ engelska
Settlementföreningen Rovalan Setlementti ry/MoniNet
värme
Äldre människor erbjuds boendeservice anordnad av Mellersta Österbottens social- och hälsovårdssamkommun Soite samt privata servicebostäder.
Sociala förmåner
Gör ditt eget videoklipp med rubriken ”Min Infobank – fem tips för dig som flyttar till Finland”.
Mer information om den ortodoxa församlingens verksamhet i Karleby finns på Vasa ortodoxa församlings webbplats.
Ansöka om medborgarskap
Information om rätten till arbetsintygfinska _ svenska _ engelska
Rättshjälpsbyråerna ger personer som är bosatta i Finland expertråd i skötseln av juridiska ärenden.
Barnet har rätt att ha kontakt med båda sina föräldrar efter skilsmässan.
Din arbetsgivare borde betala ut lönen till ditt bankkonto.
En minderårig patients åsikt beaktas när barnet är tillräckligt utvecklat för att uttrycka sin åsikt.
Läs mer på FPA:s webbplats.
Kontaktuppgifter till arbetarskyddsmyndigheternafinska _ svenska _ engelska
På InfoFinlands sida Städer hittar du information om de lokala tjänsterna i InfoFinlands medlemskommuner.
om du betalar skatt i ett annat land än Finland, din adress i det landet
Du kan börja jobba direkt när du har kommit till landet.
En sambo kan få jämkning om han eller hon till exempel genom arbete hjälpt den andra sambon att utöka sin egendom och för att det därför skulle vara orättvist att fördela egendomen enbart baserat på ägarskapet.
Boenderådgivningfinska
De bör i äktenskapet visa varandra förtroende och i samråd verka för familjens bästa.
Arbete och företagande i Finland
på ryska: 0295 020 715
efterfrågan eller säsongtopp
Innan du skaffar dig ett personligt kort ska du registrera dig som invånare i någon av kommunerna inom HRT-området.
Vid behov skriver hälsostationsläkaren en remiss till en specialist.
På rådgivningen (äitiysneuvola) följer man moderns, barnets och hela familjens välmående under graviditeten.
Omatila
familjeband
För att få rehabiliteringspenning måste du också få ett rehabiliteringsbeslut (kuntoutuspäätös) till exempel från FPA eller företagshälsovården.
Om du vill arbeta inom den offentliga förvaltningen behöver du vanligtvis ett intyg över dina kunskaper i finska eller svenska.
Du får personbeteckningen på magistraten (maistraatti) eller skattebyrån (verotoimisto).
Med hjälp av skattenumret kontrolleras, att alla arbetstagare finns i Skatteförvaltningens register.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Offentliga arbets- och näringstjänsterfinska _ svenska _ engelska
De synskadades bibliotekfinska _ svenska _ engelska
Brandsäkerhet i höghusfinska _ svenska _ engelska
ta hänsyn till arbetsgivarens intresse.
1860 Finland inför en egen valuta, mark
Att få ett förhandsmeddelande om reparationer.
Kriscentret vid Lapplands mödra- och skyddshemfinska _ svenska _ engelska
I Finland kan också två män eller två kvinnor gifta sig med varandra.
Du kan ansöka om ett banklån för detta.
Gymnasium
Den anställda på apoteket berättar för kunden om det finns ett billigare alternativ.
Läs mer på InfoFinlands sida Ekonomiska problem.
Med barnets underhållsbehov avses det penningbelopp som försörjningen av barnet kostar varje månad.
Tyska trupper som kom till Finland erövrade Helsingfors till de vita i april.
Att förlänga uppehållstillståndetfinska _ svenska _ engelska
Brand eller vattenskada
Makarna ska ingå ett avtal om barnens boende, umgängesrätt och underhållsbidrag.
EU-medborgare som har hemort i Finland kan rösta i Europaparlamentsvalet om de har anmält sig till rösträttsregistret (äänioikeusrekisteri).
För vem är yrkesinriktad arbetskraftsutbildning avsedd?
Läs mer om fastställande av faderskap vid punkten Erkännande av faderskap på den här sidan.
Anmälan till arbets- och näringsbyrån finska _ svenska
Vid servicerådgivningen får du råd och handledning utan tidsbeställning.
linkkiStiftelsetjänst:
Barn får inte l ängre cykla på trottoaren.
Man kan ansöka om Esbotillägget om en förälder tar hand om familjens alla barn under skolåldern i hemmet.
Behöver du en tolk eller översättare?
Övergången till den vanliga undervisningen sker steg för steg enligt elevens förutsättningar.
du har ett giltigt uppehållstillstånd eller uppehållskort eller att din uppehållsrätt är registrerad,
Ainonkatu 1, vån. 2
Information om gymnasieutbildningfinska _ svenska
Barnet måste ha en vårdnadshavare
De bostadslösas servicecenter på Sanduddsgatan har öppet dygnet runt varje dag.
Lönen som du får för ditt arbete kan minska ditt studiestöd.
Om personer som är bosatta i Finland antecknas grundläggande uppgifter i befolkningsdatasystemet.
Du kan boka tid för en undersökning på din egen hälsostation (terveysasema), hos en gynekolog eller på en privat barnlöshetsklinik (lapsettomuusklinikka).
Finländarna rör sig mycket till sjöss.
Enligt Finlands lag är kroppsaga mot barn förbjudet och den kan ha straffpåföljd.
Upphovsrätten till verket förblir i upphovsmannens ägo.
Lapplands läroavtalscenter ordnar läroavtalsutbildning enligt lagen om yrkesutbildning och lagen om yrkesinriktad vuxenutbildning samt stödtjänster för arbetslivet och regionutvecklingen.
Om du har flera arbetsgivare ska du förete ditt skattekort till dem alla.
Du är underhyresgäst också när du hyrt endast en del av en bostad och bostadsägaren själv bor i samma bostad.
Så här skriver du en jobbansökan och ett CVfinska _ svenska _ engelska
Man kan även studera språk.
Arbetsuppgifterna
På arbetsplatserna ska det finnas tillräckligt många personer med kunskaper i första hjälpen, första hjälpen-utrustning samt instruktioner för olycksfall.
Utbildning
Om du vill kan du skriva några ämnen på hösten och resten på våren.
Tfn 0800 414 004, tis. och ons. kl. 9–11 och 12–15
Störst är bristen på små bostäder.
linkki4V:
Tukinainen
ett annat Schengen-land begär att Finland återkallar ditt uppehållstillstånd.
Jämställdhet (tasa-arvo) mellan könen
Man kan vanligen inte få uppehållstillstånd på grund av sällskapande.
Ni kan även tillsammans besluta vem av er som tillsvidare ska bo kvar i det gemensamma hemmet.
Privat dagvårdfinska _ svenska _ engelska
Jag har inte råd att betala hyran.
du har uppgett felaktiga uppgifter i din ansökan om tillstånd
Om ditt hem är till exempel 65 kvadratmeter stort behöver du två brandvarnare.
Om bostaden har oljevärme eller elvärme, ska avgiften ibland betalas separat.
Finlands nationalspråk är finska och svenska (cirka fem procent av finländarna har svenska som modersmål).
Information om nya kurser och ansökan till kurserna finns på öppna universitetets webbplats.
Du kan be undervisningsväsendet om mer information om tjänster som skolan erbjuder.
Du kan inte registrera dig som invånare i Finland eller ansöka om registrering av uppehållsrätten när du är i landet som jobbsökande.
Vid Karleby universitetscenter Chydenius kan man avlägga såväl högre högskoleexamen som doktorsexamen.
När du är säker på att du vill och kan köpa en bostad kan du göra ett köpeanbud på bostaden.
Lär mer på InfoFinlands sida Registrering som invånare.
Detta beror dock på vilket land du kommer ifrån.
Information om spelproblemfinska _ svenska _ engelska _ ryska
Jag är dessutom rädd att jag kommer att förlora mitt uppehållstillstånd.
Navigatorn finska
Information om tuberkulosfinska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska _ bosniska _ rumänska _ swahili
Ett förmånligare alternativ till hotell är att övernatta på ett vandrarhem, men i dessa är servicenivån inte lika hög och man har inte alltid möjlighet att få eget rum.
Social-, hälso- och idrottsområdet (barnmorska, fysioterapeut, sjuksköterska)
Hur får man en delägarbostad?
linkkiPatent- och registerstyrelsen:
Du kan ringa till riksomfattande servicenummer om du behöver hjälp med att använda e-tjänsterna eller mer information om TE-byråns tjänster.
Också familjemedlemmar kan ringa eller besöka A-kliniken.
Vilka är dina styrkor?
Magistratens kontaktuppgifter och närmare anvisningar hittar du på magistratens webbplats.
Det lönar sig att söka efter en bostad på ett stort område.
Om din anställning har varat över en månad före insjuknandet betalar din arbetsgivare full lön för självrisktiden.
Alla har rätt till borgerlig vigsel, även de som tillhör ett trossamfund.
När barnet föds måste man registrera dess modersmål.
Föräldrarna kan också välja en annan skola än närskolan.
I Fpa:s beslut anges i detalj vilka omständigheter som bör anmälas.
Vardera maken ska efter förmåga bidra till familjens gemensamma hushåll och makarnas underhåll.
linkkiEira vuxengymnasium:
Flyktinghjälpens regionkontorfinska
FPA kan på din begäran föra över din ansökan om kompletterande och förebyggande utkomststöd till kommunen för behandling.
Huvudregeln är att om du bor stadigvarande i Finland, kan du få FPA:s förmåner.
linkkiFörbundet för ungdomsbostäder:
Om du säger upp bostaden den 2 juni, börjar uppsägningstiden den 30 juni och den varar en månad.
Om du reser kan myndigheterna besluta att din ansökan inte längre gäller.
linkkiAlzheimer Centralförbundet:
Maria Akademi
Som fristående examen (näyttötutkinto) (vuxenstuderande)
Helsingfors stad
InfoFinlands sidor Arbete och entreprenörskap innehåller mer information för arbetstagare och företagare.
Till din ansökan ska du bifoga:
Information om arvsskattfinska _ svenska _ engelska
Cykelkartorna är kostnadsfria.
Inledande kartläggning och integrationsplanfinska _ svenska _ engelska
linkkiAvara:
Ofta måste de som arbetar i Finland betalar skatt på sin lön i Finland.
Ärlighet och punktlighet
På FPA:s webbplats finns information om i vilka fall du kan få FPA:s pensioner utomlands.
För barn som nyligen invandrat ordnas förberedande undervisning inför grundskolan som vanligtvis pågår i ett år.
Du kan fritt välja vilken TE-byrå du besöker.
Hämta ett skattekort på den närmaste skattebyrån och lämna kortet till din arbetsgivare.
Länsi-Vantaan A-klinikka
På den här sidan hittar du information om ärenden som du måste sköta då du vill ingå äktenskap i Finland.
Intervjuerna görs i de länder där flyktingarna vistas, vanligen i flyktingläger eller i UNHCR:s lokaler.
Om det finns en vattenmätare i bostaden, fastställs vattenavgiften enligt vattenkonsumtionen.
Anmälan till språkkurserna görs vanligtvis ungefär 2–8 veckor före kursstart.
åklagarväsendet,
Dessutom måste minst två vittnen vara närvarande.
Man kan ansöka om stödet vid socialbyrån i den egna kommunen.
ådgivningarna erbjuder tjänster för gravida och barn under skolåldern.
varför du kommer till Finland (t.ex. arbete, studier)
Rådgivning om utkomstskydd för arbetslösafinska _ svenska _ engelska _ ryska
Referenser – Du kan lägga till namnen på personer som har lovat att rekommendera dig för arbetsuppgiften.
I Helsingfors trafikerar tåg, bussar, spårvagnar, metron och Sveaborgsfärjorna.
Om du vill ha en bostadsrättsbostad, hämta först ett könummer på kommunens bostadsbyrå.
Dessa telefontjänster upprätthålls av olika myndigheter och organisationer.
Också andra EU-länders medborgare som registrerat sig till rösträttsregistret i Finland har rösträtt vid Europaparlamentsval.
När ni skiljer er kan ni på förhand komma överens om hur ofta barnet kan träffa den förälder som bor på ett annat ställe.
Läs mer på InfoFinlands sida Arbetsintyg.
Patientens rättigheter
Läs mer: Gymnasium
du utvisas från Finland
linkkiUnicef:
Vid Väestöliitto får du även rådgivning på telefon eller via e-post när du behöver råd om fostran av barn eller relationerna i familjen.
Midsommar firas i slutet av juni.
Adress: Anttigatan 1, 2. våningen
grunden för de tidigare uppehållstillstånden fortfarande existerar
Du ska alltid ha ett visum när du kommer till Finland eller något annat land i Schengenområdet.
Korsholmsesplanaden 45
När uppsägningstiden har löpt ut kan hyresvärden inte kräva dig på hyra.
I skolan ges eventuellt också tilläggsundervisning, på så kallade tionde klasser (kymppiluokka).
Registreringsintyg över uppehållsrätt för EU-medborgare (om du är EU-medborgare och din uppehållsrätt måste registreras)
Läraren kan ge barnet kortvarig stödundervisning.
Om du är asylsökande i Finland eller offer för människohandel, har du rätt att få stöd för frivillig återresa (vapaaehtoisen paluun tuki), om du beslutar att återvända till ditt hemland.
Om du är intresserad av en bostad ska du kontakta något av de företag som tillhandahåller bostadsrättsbostäder:
Det uppsökande ungdomsarbetet hjälper unga i åldern 15–28 år hitta rätt tjänster till stöd för utbildning, arbete och utkomst.
Barnet lär sig även sociala färdigheter.
Läkaren kan vid behov skriva en remiss till en specialist på urologiska polikliniken.
Ibland kan arbetsgivaren också hjälpa dig med praktiska ärenden, t.ex. leta efter en bostad åt dig.
barn eller andra familjemedlemmar i Finland
1991 Den hårdaste ekonomiska krisen under
Stadsmuseetfinska _ svenska _ engelska
stöd, som man kan få när man är sjuk
Små smärtor hör till en normal graviditet när livmodern växer.
När du sköter ärenden med myndigheter, kom alltid ihåg att bekräfta tolksbehovet.
linkkiPolli.fi:
Barnet lär sig bland annat sociala färdigheter, att göra saker med händerna och olika kunskaper.
Hjälp med missbruksproblemfinska _ svenska _ engelska
Mer information om hur familjemedlemmar kan få uppehållstillstånd finns på InfoFinlands sidor Uppehållstillstånd för make eller maka, Uppehållstillstånd för barn eller förälder, Uppehållstillstånd för övriga anhöriga.
Ring inte nödnumret om situationen inte är akut.
Uppehållstillstånd eller registrering av uppehållsrätt?
Yrkesbarometern finska _ svenska _ engelska
Fråga myndigheten på förhand.
Syftet med familjepensionen är att trygga de efterlevandes utkomst.
bostadsbidraget
Förberedande undervisning tillhandahålls för invandrarbarn som inte har tillräckliga kunskaper i finska för att klara sig i förskoleundervisningen.
Utländsk yrkesexamen
Tfn 050 325 7173 (ryska, engelska)
Karleby evangelisk-lutherska församlings invandrararbetefinska _ svenska _ engelska _ ryska
Om du är under 30 år, kan du få råd och handledning via tjänsten Navigatorn.
Vårdbehovet bedöms ofta på telefon.
Inkomstregistret är en databas dit arbetsgivarna anmäler lönerna som de utbetalat till sina anställda.
Rådgivningen vid Ungdomsgården Vinge ger aktuell information om bl.a. internationalisering, studier, arbetsliv, hälsa, hobbyverksamhet och boende.
Om du behöver psykisk hjälp eller stöd, ska du kontakta din hälsostation (terveysasema).
Möblerade bostäderfinska _ engelska
Vuxensocialarbetefinska
Du kan be om råd gällande ansökan om utkomststöd via den centraliserade telefontjänsten tfn (09) 8392 1119.
När barnet fyller två år kan du inte längre använda dina faderskapspenningdagar även om sådana finns kvar.
Inom parentes anges exempel på yrken som du studera till i olika studieområden:
På en privat läkarstation måste du betala samtliga kostnader själv.
Gemensam vårdnad förutsätter att barnets föräldrar klarar av att tillsammans agera för barnets bästa.
Museerfinska _ engelska
Om det inte är fråga om ett allvarligt brott, kan du även göra brottsanmälan elektroniskt via polisens webbplats.
Tillståndsärenden
I Helsingfors finns många teatrar.
Finska medborgare som är bosatta utomlands kan också skicka vigselhandlingarna till den lokala finska beskickningen som skickar handlingarna till magistraten i Finland.
Arbetsmarknadsstödet är behovsprövat.
På MoniNets webbplats finns en studiemiljö för finska språket där du kan studera finska på egen hand.
Läs mer: Barns och ungas problem.
Du kan själv bestämma när och hur ofta du vill vara med i verksamheten.
Var särskilt försiktig om du lagar mat på natten.
Om allt är väl i övrigt kan operationen planeras i förväg.
När du kommer till Finland för att studera beror behovet av uppehållstillstånd på ditt medborgarskap.
Om du har ekonomiska problem kan du fråga om råd hos en socialarbetare i din hemkommun eller hos FPA.I vissa situationer har du rätt till utkomststöd.
Utbudet kompletteras av språk- och metodstudier.
Du kan straffas för att ha missbrukat nödnumret.
Om ditt barn plötsligt blir sjukt, ta kontakt med din hälsostation.
Fråga mer om utbudet och priserna direkt på idrottscentret.
Hobbyer för barn och unga
Inkasso
Kostnadsfri rådgivning för invandrare i frågor som rör familjens välbefinnande eller fostran av barn.
Karleby är även en betydande handelsstad.
linkkiHelsingfors och Nylands sjukvårdsdistrikt:
linkkiGuide till volontärarbete:
När du ansöker om vårdplats ska du fylla i en ansökningsblankett.
Helsingfors-info är ett rådgivningsställe där du kan fråga om aktuell information om Helsingfors, stadens tjänster, boendemöjligheter, arbete och studier.
Om du behöver akut vård samma dag, ska du ringa hälsostationen direkt då den öppnar.
Det är också bra att gå igenom bostaden och eventuella fel i bostaden med dess ägare eller hens representant.
När du bokar tid till hälsovårdstjänster kan du fråga om möjligheten att använda en tolk (tulkki) om du inte behärskar dessa språk.
Tfn 050 312 4372
Du ska ringa nödnumret endast i brådskande fall där livet, hälsan, egendomen eller miljön är i fara.
Medborgare från övriga länder måste anmäla sig personligen på TE-byrån.
Beakta att om du delar bostad med till exempel en vän och ni har ett gemensamt hyresavtal så anses ni höra till samma hushåll.
Läs mer: Tillfälligt boende.
Niande hör hemma endast i mycket formella situationer.
Företagsrådgivning fås på finska och svenska och åtminstone i de större städerna även på engelska.
På arbetspensionsutdraget finns en uppskattning av din intjänade pension.
från något annat land.
På magistraten ska du visa upp originalhandlingen eller en vidimerad kopia av den.
Uppehållstillstånd för uppstartsföretagare
Gymnasium
Höst
Lekparker och klubbar
Ett andelslag är ett företag som ägs av medlemmarna.
Familjerådgivningsbyråerna är i synnerhet avsedda för familjer med barn.
Bilagor till ansökningen ska tillhandahållas då bostad erbjuds, men kan även lämnas in tidigare.
Endast dessa familjemedlemmar kan få uppehållstillstånd på grund av familjeband.
I kollektivtrafiken kan du betala med kontanter eller resekort.
på svenska 0295 020 501
Var får jag hjälp och råd i boendefrågor?
Utlänningar som är bosatta i Finland har nästan samma rättigheter och skyldigheter som finska medborgare.
linkkiApotekareförbundet:
En ensamstående förälder fattar på egen hand alla beslut som rör barnet.
Barnet måste vara under 18 år gammalt och ogift den dag då beslutet om uppehållstillstånd fattas.
Väntetiden för dessa bostäder kan dock vara lång och endast en liten del av de sökande får en bostad.
Mer information om rätten till hemkommun finns på InfoFinlands sida Hemkommun i Finland.
Prepaid-kortet är i förväg laddat med en summa som man sedan kan ringa för.
På utrikesministeriets webbplats eller vid den närmast belägna finländska beskickningen kan du kontrollera om du behöver ett visum i Schengenområdet.
Studentexamen
Den evangelisk-lutherska kyrkan har sex finskspråkiga församlingar och en svenskspråkig församling i Vanda.
Äktenskap som ingåtts utomlands ska registreras i magistraten
Barn och ungdomar kan till exempel ha idrott, dans, musik, bildkonst eller teater som hobby.
Vid Karleby centrum finns en av landets mest omfattande historiska trästadshelheter.
Om du inte företer skattekortet till din arbetsgivare, innehåller arbetsgivaren en skatt på 60 % på din lön.
Den underlättar undersökningarna under graviditeten.
Ledande socialarbetare 016-322 3087, 040-731 2557
På mödrahemmet får du hjälp med föräldraskapet och livskompetensen.
Det är bäst att göra uppsägningen skriftligt.
Beslut om efternamn
Rovaniemi stad/idrottstjänster linkkiRovaniemi stad/idrottstjänster:
linkkiEuropass.eu:
Du kan idka många slags motion på olika håll i Helsingfors.
Information om ekonominfinska _ svenska _ engelska
Information om hemvårdsstödets kommuntilläggfinska _ svenska _ engelska
hjälper finska medborgare som råkat ut för en nödsituation utomlands
På ungdomsgårdarna ordnas också ledd verksamhet.
Läs jobbannonsen noga
Hälsotjänsterna i Helsingfors
Mer information om övriga beskattningsärenden: linkkiVerohallinto:
att kontrollera sina egna uppgifter i patientjournalen och rätta till dem
På vändagen den 14 februari kan man minnas sina vänner till exempel med blommor eller ett kort.
När du lämnar in en bostadsansökan kan du behöva också andra dokument som bilagor till ansökan.
När du bor i Finland stadigvarande, skickar Skatteförvaltningen ett nytt skattekort till dig varje år i januari.
Trettondagen den 6 januari är julens sista dag.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet
Att överklaga ett beslut om uppehållstillstånd
När ni överväger skilsmässa och behöver hjälp med att komma överens om saker och ting, kan ni ansöka om medling i familjefrågor (perheasioiden sovittelu).
Om en granne ofta bryter mot ordningsreglerna på ett allvarligt sätt, ska du först ta upp saken med grannen.
finansieringsvederlag (rahoitusvastike), om bostadsaktiebolaget har skulder
När du är sjuk
Du kan rådfråga om sådant som rör företagets verksamhet eller utveckling av företaget hos företagsrådgivningen.
Också papperslösa och asylsökande har rätt att få behandling för könssjukdomar.
linkkiEvangelisk-lutherska kyrkan i Finland:
Du kan söka dessa företag på till exempel internet.
linkkiFinlands röda kors:
I tjänsterna kan du söka information om lediga jobb och bygga upp fackliga nätverk.
På webbplatsen för Informationscentralen för teater i Finland kan du söka teatrar på olika orter på finska.
Läs mer: Brott
Läs mer på InfoFinlands sida Studier som hobby.
Diskriminering på grund av kön är förbjudet.
Du kan söka privata hyresbostäder på internet och i lokaltidningar.
Vid akuta och livshotande sjukfall kan du tillkalla ambulans genom att ringa numret 112.
Anmälan till skolanfinska _ svenska _ engelska
När du anmäler dig till skolan, kan du samtidigt anmäla dig till hemspråksundervisning och undervisning i din egen religion.
linkkiFörbundet för personaltjänsteföretag:
Läs om villkoren för familjeförmånerna på InfoFinlands sida Stöd efter barnets födelse och Stöd för vård av barn i hemmet.
Lapplands rådgivnings- och informationsservice för ungafinska
Du kan få startpenning om
Innan du startar företagsverksamheten, kontrollera om du behöver tillstånd för verksamheten eller om du måste anmäla verksamheten till en myndighet.
Då måste även de arbetsgivare som inte hör till arbetsgivarförbundet följa avtalet med sina anställda.
Du kan boka tid på rådgivningsbyrån via din hälsostation.
Läs mer: Andra studiemöjligheter
Om du har hemkommun i Finland kan du ansöka om partiell vårdpenning hos FPA för hemvård av barn under tre år eller skolbarn i årskurserna 1 eller 2.
Då läggs vanligtvis en liten förseningsavgift på räkningen.
I länder där Finland inte har en beskickning kan något annat land representera Finland i visumärenden.
om du vill studera som hobby
Du kan även få rabatt på exempelvis olika former av motion och kultur.
linkkiFinlands advokatförbund:
linkkiNödcentralsverket:
Finlands historia
Du kan använda webbtjänsten, om du har finländska nätbankskoder eller ett mobilcertifikat.
Man har hittat upp till 7 000 år gamla lämningar efter bosättning.
Under dagen får barnet en gratis måltid.
Du kan också ta ut alla 54 dagar av din faderskapsledighet vid olika tider med modern.
Den första snön kommer vanligen i oktober eller november.
Kontaktuppgifterna till invandrarbyrån i Rovaniemi är:
TE-byrån tillhandahåller tjänster som stöder utvecklingen av affärsverksamheten.
Hälsan
Erkännande och motsvarighet av examen
På 1200-talet flyttade många emigranter från Sverige till Esbo.
Vanda är en av de fyra kommunerna i huvudstadsregionen.
Information om val av kvotflyktingarfinska _ svenska _ engelska
Även om du inte använder bastun får du aldrig placera något på bastuugnen, eftersom detta kan orsaka en brand.
Arbetsgivaren har rätt att kräva ett läkarintyg för den tid då du är sjuk.
Praktik i Finlandfinska _ svenska _ engelska
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
störa eller skada fågelbon eller fågelungar
mån–tis kl. 13–21
Instruktionsfilmer om att rösta
Om du inte har pengar till bostadsrättsavgiften kan du ansöka om lån från banken.
Om du har problem i parförhållandet kan du söka hjälp vid till exempel familjerådgivningen eller hälsovårdscentralen i din hemkommun.
Ansök om tillståndet innan ditt uppehållstillstånd för studerande löper ut.
Fritidsintressen, förtroendeuppdrag
Om du vill ansöka om en hyresbostad, fyll i en ansökningsblankett för hyresbostad på Espoon Asunnot Oy:s webbplats.
Om din arbetsgivare inte betalar dig lön för den tid som du använder för teoretiska studier har du möjligtvis rätt att ansöka om dagpenning, reseersättning och familjebidrag om du omfattas av Den sociala tryggheten i Finland.
Rättshjälpfinska _ svenska _ engelska _ ryska _ arabiska
Ullavavägen 701
Man kan även köpa gymnasieböckerna begagnade.
Tandklinikernas tidsbeställning
Det är bra att ta hjälp av en jurist när du skriver ditt testamente för att det ska vara lagligt.
Ett äktenskap som ingåtts utomlands är officiellt i Finland först när det har registrerats i befolkningsdatasystemet i Finland.
Första hjälpen-anvisningar vid förgiftningfinska _ svenska _ engelska
På sommaren är det ljust i Finland även på kvällen och natten, eftersom solen går ner sent och går upp tidigt.
Ta med dig följande när du besöker magistraten:
Enligt finsk lag är alla slags diskriminering på arbetsplatserna förbjuden.
Finland förlorade kriget och var därför tvunget att betala ett tungt krigsskadestånd till Sovjetunionen i form av varor.
Nära släktingar får inte gifta sig enligt Finlands lag.
Information om presidentens uppgifterfinska _ svenska _ engelska
De ungas skyddshusfinska
Du måste dock göra en tullanmälan på flyttsakerna till de finländska tullmyndigheterna.
linkkiNyföretagarcentralerna i Finland:
Om någon upprepade gånger hotar eller trakasserar dig och du vill ha skydd, kan du ansöka om besöksförbud (lähestymiskielto) för denna person.
Om du kommer till Finland som arbetstagare någon annanstans ifrån än ett EU-land, ett EES-land eller Schweiz påverkas din sociala trygghet av följande faktorer:
FPA skickar kortet hem efter att barnet har fått en personbeteckning och ett namn.
Om du har hemkommun (kotikunta) i Finland har du rätt att utnyttja de offentliga hälsovårdstjänsterna.
Beskattningen när du börjar arbeta i Finland
Exempel:
Socialrådgivningenfinska _ svenska _ engelska
Information om finska språketengelska
Du kan använda det till exempel när du ska öppna ett bankkonto i Finland.
För att få uppehållstillstånd för uppstartsföretagare måste du ha en konkret affärsverksamhetsplan.
Julklapparna delas oftast ut på julafton.
Kontaktuppgifterna till barnatillsyningsmännen finns på Esbo stads webbplats.
Om du vill kan du ta med dig din partner till läkarmottagningen.
Om du flyttar till Finland från ett annat EU-land behöver du vanligen inte betala tull eller mervärdesskatt på dina flyttsaker, d.v.s. de personliga föremål som du tar med dig.
I Vanda beslutas ärenden av stadsfullmäktige (kaupunginvaltuusto).
Finland har två officiella språk, finska och svenska.
De centrala stegen när man startar ett företag:
Under VALMA-utbildningen kan du även förbättra dina språkkunskaper i finska.
Läs mer på InfoFinlands sida Hyresbostad.
_ holländska _ kroatiska _ rumänska _ ungerska _ italienska
Var kan jag läsa svenska?
Boendetjänsterfinska _ svenska
Naturbruk- och miljöområdet (skogsbruksingenjör, landskapsplanerare)
Adress: Porkalagatan 13 G, vån 2
På en privat läkarstation måste du betala samtliga kostnader själv.
linkkiFinlands översättar- och tolkförbund:
I ett höghus finns ordningsreglerna oftast i trapphuset.
Om du redan har uppehållstillstånd i Finland utifrån en annan grund, till exempel familjeband, kan du ha rätt att arbeta i Finland.
Du behöver inget uppehållstillstånd i Finland om du har ett uppehållstillstånd som beviljats i ett annat EU-land och om du studerar vid en högskola.
Efterforskning av anhörigafinska _ svenska _ engelska _ ryska _ somaliska _ spanska _ persiska _ arabiska _ portugisiska
Hjälp vid våld
Mer information finns på magistratens webbplats.
Tfn (09) 50 561 (växel)
via Inkomstregistrets ärendehantering, till vilken man får tillträde med webbankkoder eller andra medel för elektronisk identifiering.
Efter att en person dött kan dennes änka eller änkling och barn få familjepension (perhe-eläke).
Till långtidssjuka eller handikappade kan FPA betala ut vårdbidrag för pensionstagare.
Ansökan om dagvårdsplatsfinska _ engelska
Enligt lagen måste den som säljer bostaden berätta om de fel som han/hon känner till innan försäljningen av bostaden.
Arbetsgivaren är skyldig att trygga de anställdas säkerhet.
Tillfällig vård av barn
Anmäl ändringar till Fpa
Omskärelse får endast göras av en legitimerad läkare.
Filmklipp om tjänster inom mental hälsafinska _ engelska _ somaliska _ arabiska
Telefon: (06) 8287 750
Telefon: 040 8065 169, 040 8065 168
Entresse bibliotek, Iso Omena bibliotek, Stensvik bibliotek, Sello bibliotek och Hagalunds bibliotek.
Studierna kan även vara tilläggsutbildning eller påbyggnadsutbildning alternativt studier vid universitet eller yrkeshögskola.
linkkiVästra Nylands tingsrätt:
Det kan också finnas dolda fel i bostaden.
Polisen
Språkexamenstillfället pågår 3–6 timmar.
För att kunna bo kvar i Finland ska du ha ett jobb eller någon av de ovan nämnda anledningarna samt tillräckliga medel för din försörjning i Finland.
Information om påverkanfinska _ svenska _ engelska
linkkiRättshjälpsbyrå:
Om du är medborgare i något av de nordiska länderna, ett EU-land, ett EES-land eller i Schweiz och kommer till Finland för att studera, måste du registrera din uppehållsrätt.
Grundläggande undervisning
Kristliga folkhögskolanfinska _ engelska
Stadens hyresbostäder är förmånligare än bostäder som hyrs ut av företag och privatpersoner.
De evangelisk-lutherska församlingarna i Karlebynejden erbjuder även sorggrupper.
Människohandel är ett brott i Finland.
Läs mer: Museer.
Du kan ladda ned appen i applikationsbutiken.
I Helsingfors har man nära till naturen.
Du kan ringa om du har blivit utsatt för våld i familjen, sexuellt våld eller hot om våld.
Kom överens om när du kan gå och titta på bostaden. En bostadsvisning ordnas oftast för alla intresserade på samma gång.
Kan jag bli av med uppehållsrätten?
Bekanta dig med de lokala tjänsterna på sidorna Arbete och entreprenörskap i Esbo och Arbete och entreprenörskap i Helsingfors.
Från varje valkrets väljs ett visst antal ledamöter.
Du kan fylla i ansökan på nätet eller skicka den per post till FPA.
Läs mer: Bibliotek.
Att äta på restaurang är ofta dyrare i Finland än i andra länder.
Anmälan ska göras senast fem dagar efter löneutbetalningen.
Efter hyrestiden köper du bostaden och den blir din egen.
Det är inte nödvändigtvis möjligt att sköta alla ovannämnda ärenden i alla beskickningar.
Hälsostationerna har öppet mån–fre kl. 8.00–16.00.
Förfallodagen har antecknats i hyresavtalet.
Erkännande av examen betyder ett avgörande om vilken behörighet en utländsk examen ger när man söker jobb eller studieplats i Finland.
Bostadsaktiebolaget kan inte utfärda sådana ordningsregler som står i strid med lagen eller begränsar ett normalt liv i alltför stor omfattning.
en bostadsrättsbostad
FPA (Kela) betalar ut faderskapspenning under faderskapsledigheten.
Under andra världskriget stred Finland två gånger mot Sovjetunionen på Tysklands sida.
du har fått psykiatrisk vård i minst tre månader och
Om du har avlagt grundskolans lärokurs kan du ansöka till grundskolebaserad yrkesutbildning (peruskoulupohjainen ammatillinen koulutus).
Samarbetsprojektet Verso är ett samarbete mellan Rovaniemi stad och Rovalan Setlementti ry.
På sidorna finns nyttiga praktiska råd, kontaktuppgifter och länkar till tilläggsinformation.
Föräldrar är skyldiga att ta hand om sina barn.
Avdrag vid beskattningenfinska _ svenska _ engelska
Om du arbetar, meddela arbetsgivaren skriftligt senast två månader innan du går på moderskapsledighet.
Var och en har rätt till civilvigsel, också de som tillhör något religionssamfund.
Kan man förlora sitt finska medborgarskap?
På InfoFinlands sida Diskriminering och rasism finns information om var du kan få hjälp om du har upplevt diskriminering eller blivit offer för ett rasistiskt brott.
Stadens hyresbostäderfinska _ svenska _ engelska
Mer information om museer och aktuella utställningar får du på webbplatsen museot.fi.
du är fast anställd vid ett företag som bedriver verksamhet i ett annat EU/EES-land och ska komma till Finland för att utföra tillfälligt leverans- eller underleveransarbete och ditt arbete pågår högst tre månader;
Familjemedlem till en flyktingfinska _ svenska _ engelska
Om du har ett tidsbegränsat uppehållstillstånd som beviljats på grund av familjeband, kan skilsmässan inverka på uppehållstillståndet.
Lämna eller posta blanketten till den dagvårdsenhet där du i första hand söker plats.
I befolkningsregistret registreras alla personer som bor i Finland.
Information om bouppteckningfinska _ svenska _ engelska
Hur många timmar per vecka du arbetar eller hur lång din anställning är spelar ingen roll.
finländsk härkomst
Om du röstar på förhand kan du rösta vid vilket allmänt förhandsröstningsställe som helst i Finland eller utomlands.
Alla helgons dag
Läs mer: Äldre människor.
Parlamentsledamöterna utses genom val.
Helsingforsdagen firas varje år på dagen för stadens grundande, den 12 juni.
Utländska intyg ska vanligtvis legaliseras och översättas till antingen svenska, finska eller engelska.
Serviceguide för bostadslösa i Helsingforsfinska _ engelska _ ryska _ somaliska _ persiska _ arabiska _ bulgariska
du är asylsökande i Finland och har ett giltigt resedokument som berättigar till gränsövergång.
Du kan diskutera med dem konfidentiellt.
Du kan söka till ett universitet om du har avlagt t.ex. någon av följande examina:
Också nya elever har rätt till denna stödundervisning.
Om du fortfarande inte kan återvända till arbetet kan du söka sjukdagpenning (sairauspäiväraha) hos FPA om du omfattas av den finländska sjukförsäkringen.
uppehållstillstånd och uppehållskort (om du behöver ett uppehållstillstånd i Finland)
Adressen för TE-byrån i Karleby är
Klinikens adress eller öppettider meddelas inte offentligt.
Se Fpas hemsidor för mer information.
forskare
Privata hälsovårdstjänster är avsevärt dyrare för kunden än de offentliga.
Om du behöver en specialist, ska du först boka tid hos en allmänläkare.
Arbetarskyddfinska _ svenska _ engelska
På Utbildningsstyrelsens webbplats hittar du en förteckning över de städer där examen kan avläggas.
Radio
Webbplats för Asokoditfinska
I Esbo finns både kommunala och privata daghem.
du har din egentliga bostad och ditt hem här och så länge du huvudsakligen vistas här
Du får hjälp med att göra ett slut på våldet och råd som hjälper dig att hantera situationen.
Rådgivningen för att motarbeta diskriminering betjänar per telefon.
Mer information om museerna får du från Helsingfors turistbyrå.
Om du har ett kombinerat efternamn, till exempel Virtanen-Smith, kan du under äktenskapet lämna bort ettdera namnet.
Om makarna inte bekänner sig till samma religion förrättas vigseln i magistraten och äktenskapet kan välsignas i kyrkan.
Hjälp vid hedersrelaterade konflikter
Behovsprövad rehabilitering kan till exempel omfatta
Uppehållstillstånd för återflyttarefinska _ svenska _ engelska
I Vanda kan man få förskoleundervisning på finska, svenska och engelska.
Regionförvaltningen
uppgift om de avdrag som du söker i beskattningen för innevarande år
Du kan överklaga också om du har ansökt om uppehållstillstånd utomlands.
Om ett barn eller en ung blir mobbad i skolan är det skolans skyldighet att ingripa i detta.
Med heltidsstudier avses att studierna är din huvudsyssla.
Du kan kontakta Väestöliitto när du har funderingar kring problem i parförhållandet, fostran av barn eller skilsmässa.
När du flyttar till Rovaniemi måste du registrera dig som invånare i kommunen.
Det lönar sig att jämföra olika tjänsteleverantörers priser innan man ingår ett avtal.
Företagarens sjukdagpenningfinska _ svenska _ engelska
Du kan även få en finsk personbeteckning vid:
Om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du söka dig till en privat läkarstation.
Också ett barn som föds i Finland och blir medborgare i ett EU-land, Liechtenstein eller Schweiz måste ansöka om registrering av uppehållsrätten.
Kontrollera att du har ansökt om alla sociala förmåner som du har rätt att få.
leda arbetet och ge råd och utfärda bestämmelser som ansluter till utförandet av arbetet
För att du ska kunna få en finsk personbeteckning måste dina uppgifter registreras i Finlands befolkningsdatasystem.
Om till exempel läroanstalten ordnar dig en gratis bostad och även gratis måltider behöver du ha en mindre summa i disponibla medel.
PB 8183
Varje barn och ung person har rätt att gå i skola.
linkkiHelsingfors stadsbibliotek:
Besläktade språk är till exempel norska, danska och tyska.
På andelslagets stämma har varje medlem en röst.
linkkiCentrum för grannmedling:
linkkiTTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda:
I samband med att en integrations- eller sysselsättningsplan upprättas för dig, kan du också få också en studieplats på en finskakurs reserverad eller också kan du ställas i kö för en studieplats.
Läs mer om jobbsökning i Finland på InfoFinlands sida Var hittar jag jobb?
Det kan hända att föräldrarna förväntar sig att flickor beter sig på ett annat sätt än pojkar.
linkkiÅboregionens tolkcentral:
Läs mer: Problem med uppehållstillstånd.
Kommunen ordnar regelbundna tandläkarkontroller för barn.
Via Rovanapa Oy kan du ansöka om en bostad vid Kunta-asunnot Oy. Lediga bostäder och ansökningsblanketter hittar du även på Kunta-asunnot Oy:s webbplats..
röstberättigade personer som har grundat en valmansförening.
Paret kan hålla förlovningen privat eller offentliggöra den till andra människor.
Arbetsmarknadsstödet beviljas och utbetalas av Fpa.
Ta reda på begränsningarna också om du vill beställa läkemedel till Finland per post.
Du kan studera finska eller svenska.
En sjuksköterska eller läkare svarar i telefonen.
linkkiEsbo kyrkliga samfällighet:
Du får inte heller lägga avfall från exempelvis ditt företag i sopkärlen avsedda för ditt eget hus.
Dessutom ska den ifrågavarande kommunen vara din hemkommun senast den 51:a dagen före valdagen.
Hälsostationenfinska _ svenska _ engelska
Arv vilkas värde understiger 20 000 euro är skattefria.
Innan du flyttar in som underhyresgäst ska du säkerställa att hyresgästen har rätt att ta en underhyresgäst.
Att söka till gymnasiet
Om du har avlagt en yrkesexamen utomlands kan du ansöka om ett utlåtande om det hos Utbildningsstyrelsen.
Nyföretagarcentralen Firmaxifinska
Läs mera på InfoFinlands sida Arbetsgivarens rättigheter och skyldigheter.
Jouren har öppet varje dag dygnet runt.
Du måste alltid lämna in en separat ansökan till FPA om de socialskyddsförmåner som du behöver i din livssituation.
Om du vårdar barnet i hemmet har du rätt att ta ut oavlönad vårdledighet från ditt arbete ända tills barnet fyller tre år.
När du har fått ett könummer, kan du höra dig för om lediga bostäder hos ägare och byggherrar.
linkkiBrottsofferjouren:
Du kan inte heller ansöka om privatvårdsstöd för den kommunala småbarnspedagogiken.
Bostadsaktie
Sidorna är enkla att använda med olika enheter, till exempel smarttelefonen eller surfplattan.
En person som inte kan bo på egen hand kan bo på en anstalt.
Information om Europaparlamentsvalfinska _ svenska _ engelska
rådgivning om arbetspension och om A1-intyget
Finland är en republik och medlem i Europeiska unionen (EU).
Personer som har sin hemkommun i Esbo kan få hemvårdens stödtjänster av Esbo stad, till exempel måltidstjänster eller färdtjänst.
Om du tar hand om en äldre, sjuk eller handikappad anhörig hemma så att hen ska kunna bo hemma, kan du ha rätt till stöd för närståendevård.
Läs mer: Barns och ungas problem
Fyrverkeripjäser kan köpas i affären.
Vanligen kan man få tillstånd om man är make/maka, sambo, minderårigt barn eller förälder till minderårigt barn till personen bosatt i Finland.
De samiska språken tillhör urspråken i Finland.
byta en hel enfas anslutningsledning (spänning 230 V) och stickkontakt i en elapparat, om den gamla gått sönder.
Kommunalval förrättas vart fjärde år.
I Karleby finns stadens egna daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Fpa har en telefontjänst för barnfamiljer.
Läs mer: Officiellt intyg på språkkunskaper.
Värst var depressionen i början av 1990-talet, då det fanns ett stort antal arbetslösa i Finland, många företag gick i konkurs och staten hade lite pengar.
Missbruks​problem
En rörelsehandikappad person kan inte röra sig självständigt eller utan hjälpmedel.
I Finland är det också viktigt att man håller fast vid tider.
En cykelkarta i pappersformat för Vanda kan du hämta i Vandainfo.
Du kan också lägga till ett fotografi.
linkkiDiabetesförbundet:
Delägarbostad
PB 1002, 67101 Karleby
Vad är diskriminering?
Om du inte kan komma överens om saken med säljaren, ta då kontakt med konsumentrådgivningen.
Personer ntresserad av friluftsliv bör läsa mer om allemansrätten under rubriken ”Att röra sig i naturen” i denna tjänst.
Du måste dock studera på heltid och framskrida i dina studier.
Du kan även skicka e-post.
Med arbetslöshetsförmånen understöds bara heltidsstudier.
Information om beskattningenfinska _ svenska _ engelska
Oy Hyresboende
Guiden Bli företagare i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska _ kurdiska
Patientavgifterfinska _ svenska _ engelska
Du får inte installera en diskmaskin själv, utan arbetet måste utföras av en fackman.
Grundläggande utbildning för vuxna invandrarefinska
En del flyktingar väljs utan intervju på basis av UNHCR:s dokument.
Du behöver ett bankkonto för att sköta din dagliga ekonomi.
Verksamhetsställen för handikappservicefinska _ svenska _ engelska
Du ska lämna in en redovisning, exempelvis läkarintyg eller utlåtande från familjerådgivning.
Genom testamente kan de säkerställa att en viss egendom, till exempel den gemensamma bostaden, ärvs av sambon.
Utan tidsbokning kan du besöka Kipinä på tisdagar och onsdagar kl. 12.00–18.00.
Invandrarbyrån
Därtill är det möjligt att i vissa fall få tjänster som är särskilt avsedda för äldre.
Till Finland som företagare
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Med uthyrning i andra hand avses att hyresgästen hyr ut hela bostaden till en annan person.
på finska till numret 01019 5202 må-fre kl. 9–7, på veckoslut och helger kl. 15–7
Läs mer på InfoFinlands sida Jämlikhet och jämställdhet i arbetslivet.
Om du inte hittar en förmånlig bostad där du vill bo, fundera om du kan tänka dig att bo i en mindre bostad eller längre bort från centrum.
Moderskapsledighet
Rådgivning på engelska: 0295 020 713
Arbetsavtalslagenfinska _ svenska _ engelska
Mer information om sjukdagpenningen får du på FPA:s webbplats.
linkkiForenom:
Även försäkringsbolag, banker och många privatpersoner hyr ut bostäder.
Du kan fråga din pensionsanstalt eller Pensionsskyddscentralen om råd.
Vårdnad om barn och umgängesrättfinska _ svenska
Om barnet har feber eller annars är sjukt ska det inte tas till dagvården.
Om du inte är säker på om du har rätt till hemkommun i Finland kan du kontrollera detta vid magistraten.
Rättshjälp till brottsoffer
Välj efternamnet redan när ni ansöker om prövning av hinder mot äktenskap.
Vad ska jag göra om jag inte har hemkommun i Finland?
Partiell vårdpenning betalas inte för vård av ett barn som fyllt tre men ännu inte går i skolan.
Sexuella minoriteter och könsminoriteters rättigheter
tfn 016 322 2538
Lagen om likabehandling (yhdenvertaisuuslaki) förutsätter att alla arbetssökande behandlas lika.
I vissa fall får du en tolk via myndigheten.
På deras webbplatser kan du också ladda ned företagarhandböcker åtminstone på finska och på engelska.
Barnskyddet har många slags medel som de kan använda för att hjälpa familjen.
Tfn (09) 5056 297
Delegationen för mångkulturella frågorfinska
Ortodoxa församlingenfinska _ ryska
Hur får jag ett tillfälligt uppehållstillstånd ändrat till ett kontinuerligt tillstånd?
Mental hälsa
Du kan använda mödrarådgivningstjänsterna i din hemkommun om du har hemkommun (kotikunta) i Finland.
Översättningsanvisningen är på finska.
Välja efternamn
Barnets vårdnadshavare har även rätt att få information om allt som berör barnet av myndigheter.
Om
Boende i en krissituation
Fundera också på hur du ordnar bokföringen och planerar ekonomin.
din flyktingstatus i Finland har upphört eller återkallats eller det har fattats beslut om att avvisa dig.
Läs mer på InfoFinlands sida Om du blir arbetslös.
Medborgarinstituten och arbetarinstituten ordnar finskakurser för invandrare.
Från fackförbund får du mer information om lönenivån i olika branscher.
Kurser hålls på finska, engelska och ryska.
forskaruppdrag
Barns hälsa
Företagarnas stödnät (Yrittäjän tukiverkko) är en gratis webbtjänst som Företagarna i Finland upprätthåller. Tjänsten innehåller mycket nyttig information för företagare.
språk
Läraren lär känna eleverna bra och kan utveckla undervisningen så att den passar dem.
Språkkurserna är ofta fullsatta.
Kontakta rådgivningsbyrån (neuvola) när du upptäcker att du är gravid.
I det finländska samhället är alla jämlika och alla ska behandlas rättvist.
Storleken av försäkringspremierna och pensionen beror på hur stor förvärvsinkomst (työtulo) förtagaren har.
Kontrollera i lönespecifikationen och skattedeklarationen (veroilmoitus), att arbetsgivaren har betalat skatt på din lön.
För föreningen väljs en styrelse på föreningsmötet dit alla föreningsmedlemmar sammankallas.
Berätta på ditt sätt vad som är bra att veta när man ska flytta till Finland.
Smärtor och blödningar under graviditeten
I Finland föder kvinnorna vanligen på sjukhus.
Studerandehälsovårdfinska _ svenska
Därefter fattar Migrationsverket beslut om uppehållstillstånd.
Simpass för invandrarkvinnorfinska _ engelska
Elektronisk ansökanfinska _ svenska _ engelska
Penningunderstöd och stipendier
Du ansöker om studiepenning och statsgaranti för studielån vid FPA.
Arbets- och näringsbyrån hjälper dig i jobbsökningen.
Mer information om dessa museer finns under länkarna här intill.
Vid rådgivningarna utförs vaccinationer av barn och vuxna.
Då minns man Jesu himmelsfärd.
Om du blir bostadslös ska du kontakta socialbyrån eller socialstationen i din hemkommun.
I skyddshemmet är du i säkerhet och där finns personal på plats hela tiden.
Man kan ringa eller besöka Nupoli.
När samboförhållandet upphör delas egendomen vanligtvis så att båda parterna får sin egen egendom.
Information om tandvårdsjourenfinska _ svenska _ engelska
Information om gränssnittetfinska _ engelska
är införd i befolkningsdatasystemet
Kollektivtrafik
Hjälp för kvinnor för att sluta med våldsamt beteendefinska _ svenska _ engelska
01301 Vanda
Du får mer information om dessa standardblanketter hos myndigheterna i det land där du begär intyget.
När barnet blir sjukt ska du vid behov kontakta Grankulla hälsostation.
Basfakta
Information om tjänster som underlättar vardagen för äldre får du på InfoFinlands sida Äldre människor.
I stadsfullmäktige sitter 75 ledamöter som representerar olika politiska grupper.
Lag om hemkommunfinska _ svenska
Det är det billigaste sättet att resa.
De lär sig nya saker med lekens hjälp.
Om du är medborgare i något EU-land, Liechtenstein eller Schweiz och flyttar till Finland permanent, ska du registrera dig vid Migrationsverket och magistraten.
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en krismottagning för invandrare som bor i Helsingforsregionen.
Tandsjukdomar behandlas på bästa sätt då de upptäcks innan symptom uppkommer.
Filmerfinska
Om om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du gå till en privat tandläkare.
Tjänsten ger service på finska, svenska och engelska.
Förskoleundervisningen ges av pedagoger inom småbarnsfostran som har avlagt universitetsexamen.
Blanketter för ansökan om uppehållstillståndfinska _ svenska _ engelska
I Rovaniemi finns ungdomsgårdar i åtta olika områden: centrum, Korkalovaara, Nivavaara och Ylikylä samt byarna Muurola, Sinettä, Oikarainen och Vanttauskoski.
Tandvårdens nattjour (hammashoidon yöpäivystys) finns på Tölö sjukhus olycksfallsstation.
linkkiSeta:
linkkiEnergimarknadsverket:
Du kan hyra en bostad av privata hyresvärdar eller ansöka om en av Helsingfors stads hyresbostäder.
Studier i finska språket på Internetfinska _ engelska
Företagshälsovårdfinska _ svenska _ engelska
Socialrådgivningen (sosiaalineuvonta) ger information om utkomststöd (toimeentulotuki) och andra bidrag om du har ekonomiska problem.
I Esbo finns flera läroanstalter som ger grundundervisning i konstämnen speciellt för barn och unga.
Kvällstid och under veckoslut har hälsostationerna stängt.
Övrig undervisning i Karlebyfinska _ svenska
Information om öppna yrkeshögskolanfinska _ svenska
Serviceguide för bostadslösa i Helsingfors(pdf, 3,7 MB)finska _ engelska _ ryska _ somaliska _ persiska _ arabiska _ bulgariska
att organisera sig
Via en patientförening kan man också hitta kamratstöd.
På din egen hälsostation får du mer information om hur mentalvårdstjänsterna är ordnade i din hemkommun.
Arbets- och näringstjänsten
Ring inte nödnumret om ärendet inte är brådskande.
Om du har avlagt en examen i Finland kan du få ett tillfälligt uppehållstillstånd för arbetssökande.
Stöd för närstående till rusmedelsberoende personerfinska _ svenska
Nyår
Om du blir tvungen att betala kvarskatt, får du tillsammans med beskattningsbeslutet en bankgiroblankett.
Bostadsförmedlaren kräver att jag betalar hen för att få se bostaden.
Tjänsten kan till exempel vara att du får hjälp med att leta efter en bostad eller arbetsplats i det land dit du återvänder.
Konst Vionojafinska
Om ditt barn har en specialdiet ska du tala om det för läraren.
Stöd för lärande arrangeras i mån av möjlighet på elevens eget modersmål i skolan.
Röda Korset hjälper familjer som skilts åt vid olika katastrofer eller kriser.
Barnet eller den unga kan även delta i förberedande undervisning.
Till exempel kan mamman till ett litet barn förvärvsarbeta medan den andra föräldern stannar hemma för att ta hand om barnet.
Miehen Linja betjänar på finska, engelska, svenska, franska och grekiska.
En utredning över att du har betalat läsårsavgiften eller har ett stipendium
Största delen av finländarna bor ägarbostäder.
Hemvårdsstöd för barn och Helsingforstilläggetfinska _ svenska _ engelska
Föreningen för små familjer är en medborgarorganisation som grundats av ensamstående föräldrar och som erbjuder aktiviteter för medlemsfamiljerna.
Flyttfirmor
Hemstadsstigarfinska _ svenska _ engelska
Runebergsdagen
bilskatter
om du söker till ett magisterprogram
I detta fall står det i bolagsordningen vem som ansvarar för vad.
Om du är i akut behov av vård, ring tidsbeställningen direkt på morgonen.
Du kan även skicka in ansökan till tingsrättens kansli per post, som telegram eller via e-post.
Via TE-byrån kan du även leta en fortsättare för din företagsverksamhet eller en partner till ditt företag.
Man kan också ordna en civil begravning utan religiösa inslag.Om civil begravning får du information hos servicecentret Pro-Ceremonier (Pro-Seremoniat).
Eget initiativtagande och ansvar
Småbarnspedagogiken ordnas i daghem och familjedagvården.
Ansökan till VALMA-utbildningfinska _ svenska
Hälsovård för EU-medborgare
Uppsägning av bostad
Om du har barn och ska skilja dig tar du kontakt med barnatillsyningsmannen (lastenvalvoja) vid Vanda stad.
I Vanda kan du studera på gymnasiet (lukio) på finska, svenska eller engelska.
I tillgången till dagvårdstjänster är målet att uppfylla närserviceprincipen för varje barn.
På adressen Ilmonet.fi hittar du hela kursutbudet vid arbetar- och medborgarinstitut i huvudstadsregionen.
De rusmedels- och rökfria ungdomslokalerna erbjuder handledd verksamhet för barn i årskurserna 3–6 och unga i åldern 13–17 år i olika delar av Karleby.
Företag som har förutsättningar för lönsam verksamhet, men inte den egenfinansieringsandel eller de garantier som bankerna kräver, kan få ett lån eller borgen för ett lån vid Finnvera.
Om du arbetar permanent kan du även ansöka om uppehållstillstånd i Finland på grund av arbete.
tortyr eller någon annan behandling eller bestraffning som är omänsklig eller kränker människovärdet eller
Seure erbjuder kortvariga jobb vid Helsingfors, Vanda, Esbo och Grankulla städer.
På Vandakanalen kan du följa fullmäktiges sammanträden och få mer information om beslutsfattandet.
Kommuner, församlingar och vissa organisationer ordnar nödinkvartering.
Behöver du en jurist?
Om du bor i Finland tillfälligt, registreras ingen hemkommun för dig i Finland och du har inte samma rättigheter som de personer som bor i Finland stadigvarande.
Anteckna i affärsverksamhetsplanen också hur du tänker ordna bokföringen och ekonomiplaneringen och hur du följer upp realiseringen av dina planer.
Arbetsgivare måste också ge arbetstagaren ett nytt arbetsintyg om arbetstagarens arbetsintyg kommer bort eller förstörs.
Migrationsverket ger rådgivning angående tillstånd också per telefon.
linkkiBefolkningsförbundet:
Omskärelse och förlossning
Om det är fråga om ett allvarligt brott, kan polisen gripa eller anhålla den brottsmisstänkta.
Portugisiska
linkkiKonsumentförbundet ry:
Då kan bodelningen jämkas.
Kravet om att äktenskapet ska dömas till skilsmässa efter betänketiden görs likadant som den första ansökan.
Både arbetsgivaren och den anställda undertecknar arbetsavtalet.
Via tjänsten kan du också fråga om anvisningar för vård av sjukdomar.
yrkesinriktade grundexamen, yrkesexamen eller specialyrkesexamen
Du behöver Utbildningsstyrelsens eller någon annan myndighets beslut om erkännande av examen om du vill arbeta inom ett reglerat yrke eller en uppgift som kräver högskoleexamen på viss nivå.
Då får du en finsk personbeteckning på samma gång som du får uppehållstillståndet.
Legalisering och översättning av intyg
Skolpsykologerfinska _ svenska
Motionsplatserfinska _ svenska
Använd inte material, såsom bakgrundsmusik eller bilder, som en tredje part har upphovsrätt till.
I Grankulla tillhandahålls offentliga hälso- och sjukvårdstjänster på hälsostationen.
Om du inte har möjlighet att identifiera dig i Mina e-tjänster eller om du vill uträtta dina ärenden per telefon kan du få information, rådgivning, vägledning och stöd i användningen av nättjänsterna från den nationella telefontjänsten.
Hjälpmedel
På rådgivningen diskuteras parförhållandet och föräldraskapet samt papparollen och föräldrarnas ansvar.
Jobbsökning i Finland
Yrkesutbildning ger den studerande behörighet till ett visst yrke.
I och med produktionen av krigsskadeståndet utvecklades
Dessa examina avläggs alltid genom fristående examen.
Ett delbeslut av arbets- och näringsbyrån behövs inte för tillståndet.
Avvisning av en asylsökandefinska _ svenska _ engelska
När användaren är på en kommunsida, visas länkar till den grundläggande informationen om ämnet.
Helsinki-info betjänar på många olika språk per telefon, ansikte mot ansikte och elektroniskt.
Tjänster för företagare-Startup Kitfinska
Om du är turist i Finland och hamnar i en svår situation, ska du kontakta ditt hemlands beskickning.
Tack.
När du ansöker om uppehållstillstånd, kan du samtidigt även ansöka om en finsk personbeteckning.
Begravningsplatserfinska _ svenska
Bioavfall (biojäte)
Vid ett olycksfall i skolan får barnet första hjälpen.
Priser på icke subventionerade hyresbostäderengelska
Om du betalar för litet i skatt, blir du tvungen att betala kvarskatt.
De som är klienter vid FPA kan få utbildningsstöd under utbildningen.
Alla som vill lära sig tala finska är välkomna till caféerna.
Vår
Om du reser i hemlandet eller utomlands ska du se till att du alltid kan nås.
linkkiDiskriminerings- och jämställdhetsnämnden:
När du flyttar till Finland ska du besöka magistraten (maistraatti)på orten där du är bosatt.
Tfn (09) 839 35013
Inkomstregistret
I anmälan anges barnets närskola (lähikoulu).
linkkiFörbundet för ungdomsbostäder:
linkkiArbis:
Om din anställning varat över en månad före insjuknandet får du lönen till fullt belopp för minst den dag då du insjuknade och nio därefter följande dagar.
svara på nödcentraloperatörens frågor
Arbetsgivaren ansvarar för att alla kan arbeta tryggt.
Läs mer: Problem med uppehållstillstånd
arbetssituation
Du kan besöka Karlebynejdens Utveckling Ab om du behöver information om att grunda ett företag.
Information om integrationfinska _ svenska _ engelska
På webbplatsen för evangelisk-lutherska kyrkan i Finland hittar du information om kyrkans tjänster.
På InfoFinlands sida Komihåglista för dig som flyttar till Finland hittar du nyttig information om allt som du ska ta hand om när du flyttar till Finland.
På Seniorrådgivningen (seniorineuvonta) får du information om hobbyer och tjänster för seniorer som olika organisationer, företag och staden erbjuder.
Vad stadigvarande boende betyder definieras i lagen.
Om du är 17–64 år gammal och på grund av din livssituation inte har anmält dig som arbetslös arbetssökande kan personalen på Rovaniemi stads socialservicecenter göra en inledande kartläggning och vid behov även en integrationsplan tillsammans med dig.
Om inkomsten som man får för försäljningen av varor och tjänster är mindre än 10 000 euro per år, behöver ingen mervärdesskatt betalas på den.
Exempelvis föräldrarna har inte rätt att tvinga eller utöva påtryckning på sitt barn att gifta sig.
TE-byrån i Österbotten betjänar i Karleby, Kaustby, Jakobstad, Närpes, Kristinestad och Vasa.
Santa Sport Spafinska
Information om hemvårdens stödtjänsterfinska
Var och en har alltså rätt att bekänna och utöva sin religion.
Vårdnaden om ett barn innebär
De tysta stunderna behöver inte fyllas med prat.
I Helsingfors erbjuds tolktjänster av flera företag.
Det är även möjligt att ett existerande tillstånd upphävs.
Du får mer information i skolan.
Olika skolor
Det är viktigt att du även själv aktivt främjar din integration.
Bostadsaktiebolaget ska se till att husets konstruktioner, isolering, värmesystem, elledningar, vattenledningar och avlopp samt gårdsområden hålls i gott skick.
I dag finns det många medborgarorganisationer som specialiserat sig på att främja en viss samhällelig fråga.
Du kan komma direkt till SERI-stödcentret på egen hand, men det rekommenderas att man ringer i förväg.
Förenta nationernas flyktingorganisation UNHCR. Kvotflyktingarna väljs bland de personer som UNHCR föreslår till Finland.
Hyresvärden föreslog att vi gör ett muntligt hyresavtal.
Läs mer: Barns hälsa.
Högljutt prat kan anses vara obekvämt eller hotfullt.
Hur mycket de olika sidorna används
Vid hälsostationen får du mer information om hjälpmedlen.
Du hittar de separata ansökningarna via tjänsten Studieinfo.fi.
Hyresbostäderna är ofta dyra i huvudstadsregionen.
Dessa kan inte underskridas i arbetsavtalet.
Om du flyttar till Finland av familjeskäl omfattas du vanligen av det finländska socialskyddet.
Om du har svårt att sköta din ekonomi, betalningssvårigheter eller skulder kan du få råd av en ekonomi- och skuldrådgivare.
Målargränden 3 B
Vissa tolkcentraler håller vid behov jour på veckoslut och kvälls- och nattetid och även med kort varsel.
Vid Kronoby folkhögskola kan du studera finska och svenska på grund- och påbyggnadsnivå.
Videoklippet får inte vara kränkande, nedsättande eller diskriminerande mot kön, etniskt ursprung eller religiös övertygelse.
Medborgarrådgivningen guidar dig till den rätta tjänsten, hjälper med digital ärendehantering och besvarar allmänna frågor om de offentliga tjänsterna.
Uppsägningstiden gäller hyresavtal som gäller tillsvidare.
Du kan söka information om möten på webbplatsen på finska, engelska och svenska.
Dessutom måste dina studier:
Föreningens verksamhet
I samma val kan du rösta i endast ett EU-land.
Barnets medborgarskap påverkar inte huruvida du får stöd eller ej.
Inledande kartläggning och integrationsplan
Rådgivningarnas telefontjänst
Hälsovårdaren på rådgivningsbyrån frågar om du har blivit utsatt för könsstympning.
Läs mer: Bostadsrättsbostad.
Stäng alltid av en elektrisk bastuugn efter användning.
Stäng alltid av en elektrisk bastuugn efter användning.
Regnbågsfamiljer
Förskoleundervisning i Helsingforsfinska _ svenska _ engelska
Information på webben
Anvisningar om ansökning och närmare information om utbildningsprogrammen finns på högskolornas egna webbplatser.
linkkiBab.la:
Viktiga händelser
Om någon annan hälsovårdsenhet behöver dina uppgifter, ombeds du ge ditt medgivande för överlåtelse av dessa.
De flesta är finskspråkiga.
Begravning
Registreringen hos Migrationsverket är inte samma sak som registreringen av din bosättningsort i befolkningsdatasystemet (väestötietojärjestelmä) vid magistraten (maistraatti).
Du hittar information om körkort på polisens och Trafiksäkerhetsverkets (Liikenteen turvallisuusvirasto) webbplatser.
Du får en personbeteckning av Migrationsverket när du beviljas uppehållstillstånd i Finland eller när din uppehållsrätt för EU-medborgare registreras.
Företagsrådgivningfinska _ engelska
Åldringar som dagligen behöver utomstående stöd och hjälp har rätt till serviceboende.
Diu kan boka en tid genom att ringa hjälptelefonen i förväg eller besöka centret.
Du får mer information på InfoFinlands sida Hälsotjänsterna i Finland och Äldre människors hälsa.
Då får du en finsk personbeteckning samtidigt som du får ditt uppehållstillstånd.
Ingående av äktenskapfinska _ svenska _ engelska
Prövning av hinder mot äktenskap
Handläggning av brottsmål i tingsrättenfinska _ svenska _ ryska _ arabiska
FPA och Skatteförvaltningen erbjuder information till utländska anställda på servicestället In To Finland i Helsingfors.
Arbets- och näringsbyrån i Esbo
Varje skola har en läkare och en hälsovårdare.
I de nordligaste delarna av Finland går det flera veckor utan att solen går upp överhuvudtaget.
Du får närmare uppgifter av parktanterna per telefon.
Information om den förberedande utbildningen får du vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning.
Pass ansöks på polisstationen.
Om du behöver juridisk hjälp, kan du kontakta Västra Nylands rättshjälpsbyrå.
söker heltidsarbete
Social-, hälso- och idrottsområdet
Information om Esbofinska _ svenska _ engelska
När du tar hand om en anhörig i hemmet
Du betalar avgiften när du lämnar in din ansökan.
Du betalar för färdtjänsten enligt kollektivtrafikens taxa.
Den inledande kartläggningen hjälper dig att hitta rätt tjänster i din hemstad.
67100 Karleby
linkkiFinlands flyktinghjälp r.f.:
Om du letar efter en viss bok, kan du också be om hjälp av personalen på biblioteket.
Mer information om hemspråksundervisning och om undervisning i elevens egen religion hittar du på stadens webbplats och hos områdeskoordinatorerna (aluekoordinaattori).
Om du vill byta efternamn ska du ansöka om namnändring hos magistraten.
Information om var din närmaste återvinningsstation (kierrätyspiste) ligger hittar du på webbplatsen kierrätys.info.
Inledande kartläggning och integrationsplan
Barnlöshet
Information om medlemskortetfinska _ svenska _ engelska _ ryska _ franska _ somaliska
I allmänhet ordnas den gemensamma ansökan i februari-mars och september-oktober.
Det andra inhemska språket (finska eller svenska)
Du får faderskapspenning även om du inte bor tillsammans med barnets mor.
Kontaktuppgifter för den grundläggande utbildningenfinska
Om du bara vill hälsa på hos din familjemedlem i Finland hittar du mer information på InfoFinlands sida Kort vistelse i Finland.
Tidsbeställning per telefon mån–ons kl. 9–10.
Huvudhälsostationens tandklinik
Om du blir sjuk och inte kan arbeta ska du utan dröjsmål meddela detta till din chef.
Tfn (09) 8789 1300
Det här kallas för förskottsinnehållning (ennakonpidätys).
Medborgarinstitutet i Rovaniemi erbjuder kurser i finska språket.
Likabehandling och förebyggande av diskriminering på arbetsplatserfinska _ svenska _ engelska
Offentliga tjänster på internetfinska _ svenska _ engelska
När du köper ett telefonabonnemang i Finland får du ett finskt telefonnummer.
I Esbo anordnas förskoleundervisningen (esiopetus) i daghemmen.
Högskolorna har vissa utbildningsprogram där undervisningen ges på engelska.
Barnatillsyningsmannen ordnar ett möte med föräldrarna.
Albertinkatu 25
Det är rekommendabelt att arbetsavtalet är skriftligt.
Före äktenskapet måste en prövning av hinder mot äktenskap (avioliiton esteiden tutkinta) göras.
Du kan också lägga till sådant kunnande som du har införskaffat till exempel i frivilligarbete, fritidsintressen eller studier.
Identifiera och dra nytta av dina nätverk.
I Mina e-tjänster på nätet kan du bl.a. ändra dina uppgifter som arbetssökande och kontrollera giltighetstiden för jobbsökningen och utlåtandet om arbetslöshetsförsäkring.
Telefon: 050 3147 464.
Du kan ansöka om uppehållstillstånd på något av följande grunder:
hur länge arbetet varar
Den ligger mitt i Esbo, 15 kilometer västerut från Helsingfors.
På många arbetsplatser vill man stödja de anställdas arbetsmotivation och -trivsel med olika rekreationsdagar och fester på arbetsplatsen. Arbetsgivaren kan också erbjuda sina anställda olika hobbymöjligheter vid sidan av arbetet.
Inkomsten beskattas utifrån företagets förmögenhet antingen som kapitalinkomst (pääomatulo) eller som förvärvsinkomst (ansiotulo).
Du kan arbeta i Finland utan uppehållstillstånd till exempel om:
På sjukhuset samtalar en skötare och en läkare med dig.
Till samma hushåll hör vanligtvis alla som stadigvarande bor i samma bostad.
Information om företagsformerfinska _ svenska _ engelska
Du har ändå själv ansvaret för att dina fakturor skickas till rätt adress och betalas i tid.
Staten
Reservera tillräckligt med tid för att hitta en bostad.
De erbjuder utbildning inom många olika branscher.
muntliga färdigheter
Privat tandvård är dyrare än offentlig tandvård.
FPA har bland annat hand om folkpensionen, barnbidrag, det grundläggande utkomstskyddet för arbetslösa, sjuk- och föräldradagpenningar, utkomststöd och rehabilitering.
Skolmaten är gratis för alla och man behöver inte ta med sig en matsäck till skolan.
I Europeiska unionens råd är regeringarna för medlemsländerna representerade.
Läs mer om dessa förmåner på InfoFinlands sida Stöd till gravida.
Rovaniemi stads idrottstjänster erbjuder personer över 27 år (inte heltidsstuderande) möjlighet till regelbunden motion i hälsomotionsgrupper.
Många kommunicerar med teckenspråk.
Lapplands landskapsbibliotek
I den finländska kulturen framhävs individualism mer än i många andra kulturer.
Läs mer om rätten till hemkommun på InfoFinlands sida Hemkommun i Finland.
Barn har rätt till att deras åsikt tas i beaktande när man fattar beslut om sådant som rör dem.
Den ligger intill Esbo och Helsingfors.
Specialister finns på vissa hälsostationer, på polikliniker och sjukhus.
Esbo är en av huvudstadsregionens fyra kommuner.
Öppna daghem (avoin päiväkoti) är avsedda för barn under skolåldern och de föräldrar och vårdare som tar hand om dem.
Du kan endast ansöka om fortsatt uppehållstillstånd i Finland.
Du hitar mer information om föreningar på InfoFinlands sida Föreningar.
Om du upplever diskriminering någon annanstans än på jobbet eller om du har upptäckt diskriminering någonstans kan du ta kontakt med diskrimineringsombudsmannen (yhdenvertaisuusvaltuutettu).
Lediga bostäder och ansökningsblanketter hittar du även på Kunta-asunnot Oy:s webbplats..
Social- och krisjouren vid Jorv sjukhus i Esbo hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation, till exempel vid våld, problem med barnen eller psykiska problem.
försvar
Mångkulturell barndagvård i Rovaniemi betyder att alla barn beaktas likvärdigt och rättvist oavsett ålder, kön eller hudfärg.
Ohjaamo-verksamheten erbjuder råd och vägledning till unga bostadslösa.
Den egentliga dagen för firandet är julafton den 24 december.
Startpunkt för unga vuxna
Barn i skolåldern går på tandläkarkontroll under skoldagen vid tandkliniken i området.
Om du inte har tillräckliga språkkunskaper eller studiefärdigheter för yrkesutbildning, kan du före yrkesutbildningen söka till utbildning som handleder för yrkesutbildning (VALMA).
Anmäl dig som arbetssökande i TE-byråns webbtjänst.
Ansökan om Schengenvisumfinska _ svenska _ engelska
Lärarna i årskurserna 7–9 har läst det ämne som de undervisar.
Om du behöver en personbeteckning för arbete, kan du få en personbeteckning även på skattebyrån.
Du kan ladda resekortet på vilket serviceställe för resekort (matkakortin latauspiste) som helst.
I många nationalparker finns forststyrelsens naturcenter där man får aktuell information om områdets natur och om hur man ska röra sig i området.
Om du behöver en tolk, ska du uppge detta när du bokar tiden.
Om barnet går i en svensk skola kan hen läsa svenska som andra språk.
Samtalet besvaras av en sjukskötare eller en läkare.
Tandvårdens nattjour (hammashoidon yöpäivystys) finns på Tölö sjukhus olycksfallsstation.
På många orter finns också andra religionssamfunds begravningsplatser.
I arbetsavtalet står det ofta hur långa pauser som ingår i arbetsdagen och tidpunkten för dessa.
Par med barn under 13 år kan vid problem i äktenskap och parförhållande få hjälp vid familjerådgivningen (perheneuvola).
Napapiirin Residuum
Du kan också lämna in en ansökan vid ett serviceställe.
Medborgarinstituten ordnar förmånlig musikundervisning.
Filmklippet ska vara 1–3 minuter långt.
På Utbildningsstyrelsens webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
Identitetskort
På många mindre orter finns det många lediga bostäder och priserna är lägre.
Öppningsoperationen kan göras före graviditeten, när graviditeten är halvvägs eller i samband med förlossningen.
Arbetarinstituten ordnar kurser också på engelska och ryska.
Flyttsaker från länder utanför EU
Fråga på mödrarådgivningen på vilket sjukhus du ska föda.
Länkar till jobbsajterfinska _ svenska _ engelska
Du kan också kontakta din egen hälsostation.
linkkiVanda arbets- och näringsbyrå:
vägra att delta i verksamhet som konkurrerar med arbetsgivaren
Du får information om modersmålsundervisningen vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning.
Jämställdhetsombudsmannen övervakar att lagen om likabehandling av män och kvinnor följs.
Försäkringsbolag i Finlandfinska
Använd spisfläkten när du lagar mat.
Den närmaste jourmottagningen finns vid Jorv sjukhus i Esbo.
Mottagning /Kelviå
att man tar hand om och beslutar om barnets angelägenheter.
skriftliga färdigheter
lärare
I en del städer måste man själv boka tid för kontrollen.
På InfoFinlands sida Komihåglista för dig som flyttar till Finland hittar du nyttig information om vilka andra saker du bör ta hand om innan du flyttar till Finland.
Justitieministeriet kan på synnerligen vägande skäl ge tillstånd till äktenskap i de två sistnämnda fallen.
Kvällstid och under veckoslut har hälsostationen stängt.
Offentliga arbets- och näringstjänsterfinska _ svenska
Nödcentralsverketfinska _ svenska _ engelska
Vissa läroanstalter ordnar yrkesinriktad arbetskraftsutbildning särskilt för invandrare.
Försäkringar
A2 – ASE 2
Man kan också söka skilsmässa utan makens eller makans samtycke.
Serviceboende kan ordnas i vanliga bostäder, i ett servicehus, i en servicebostadsgrupp eller i någon annan form.
Nätverket Vi läser tillsammans (Luetaan yhdessä-verkosto) erbjuder undervisning i läsning och det finska språket för invandrarkvinnor.
du har fått ett negativt beslut på din asylansökan
Television
Hur fort studierna framskrider beror på dig själv.
JA: metallföremål och förpackningar som till största delen utgörs av metall
Möblerade bostäderfinska _ svenska _ engelska _ ryska
Helsingfors stads bibliotek är en del av HelMet-biblioteket.
Du kan ringa jourtelefonen dygnet runt.
Vid problem som berör barn i skolåldern hjälper till exempel skolans hälsovårdare.
Den ska göras i steril miljö.
Efter cirka 1995 började en ekonomisk tillväxt i Finland, varvid det viktigaste företaget var mobiltelefontillverkaren Nokia.
När du avslutar dina studier
Kontaktuppgifterna hittar du på Vanda stads webbplats.
Tullrådgivningen betjänar på finska, svenska och engelska.
Om du kommer till Finland för att söka jobb kan du vanligtvis inte få arbetslöshetsersättning från Finland.
Inom EU (och i Schweiz, Norge, Island och Liechtenstein) måste man söka asyl i det land, till vars territorium man kommer först.
För att få utkomstskydd för arbetslösa måste du aktivt söka jobb och vara beredd att ta emot ett jobb.
Du kan skicka in en öppen ansökan eller ringa arbetsgivaren, trots att de inte har några lediga jobb just nu.
Flyktingrådgivningen ger juridisk hjälp och rådgivning för asylsökande, flyktingar och andra utlänningar.
betalat alla avgifter som överenskommits med hyresvärden.
Hemspråksundervisningfinska _ engelska
Vanligtvis delas egendomen vid skilsmässa jämnt mellan makarna.
Detta meddelas i lokaltidningarna och på stadens webbplats.
Trots att du inte har uppehållstillstånd kan du börja arbeta tre månader efter att du har lämnat in din asylansökan;
linkkiUndervisnings- och kulturministeriet:
Om en familjemedlem är våldsam eller hotar med våld, ta kontakt med Karleby mödra- och skyddshem.
Därtill ägs hyresbostäder i Vanda av många försäkringsbolag, Kuntien eläkevakuutus och Kunta-asunnot.
Ofta krävs till exempel att djuren har fått vissa vaccinationer.
Hanteringen av ansökan är avgiftsbelagd. Avgiften ska betalas då ansökan görs.
Socialjouren
Utifrån den inledande kartläggningen görs en bedömning av om det även vore bra att göra upp en integrationsplan för dig.
arbetslivet
Social- och krisjouren
Graviditetspreventionfinska _ svenska _ engelska
Avgiften måste betalas i samband med att man lämnar in sin tillståndsansökan.
Om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd (perustoimeentulotuki) hos FPA.
TE-byråns adress i Karleby
Helsingfors företagare är företagarnas intressebevakningsorganisation som erbjuder sina medlemmar till exempel utbildning, nätverk och rådgivning.
Bolaget beviljar lån och borgen åt nya företag eller företag som redan är verksamma.
Svenskan som talas i Finland är finlandssvenska.
Om du behöver hjälpmedel ska du först kontakta din egen hälsostation.
Min anställning upphör inom kort.
Juristerna svarar på dina frågor på finska och engelska.
Om du misstänker att din arbetsgivare har diskriminerat dig på grund av ditt kön kan du be jämställdhetsombudsmannen om råd och anvisningar samt hjälp med att reda ut saken.
Så gör man till exempel om du inte har ett bankkonto.
Du kan ansöka om privatvårdsstöd (yksityisen hoidon tuki), om
Idrottsklubbarfinska _ svenska
Även de anhöriga till en spelberoende person kan få hjälp.
Samfund och företag som låter bygga delägarbostäder informerar om nya och lediga bostäder.
Kom ihåg att ansöka om fortsatt uppehållstillstånd för studerande i god tid innan giltighetstiden för det första tillståndet går ut.
Omskärelse och graviditet
När en person fyller 18 år är han eller hon enligt lagen myndig.
Stöd kan beviljas för fast bostad i Finland.
I Esbo finns en delegation för mångkulturella frågor som utvecklar stadens mångkulturella politik.
Information om VALMA-utbildningarfinska _ svenska _ engelska
Uppgifter som inte kräver en viss utbildning
Vad är ett hushållfinska _ svenska _ engelska
Du hitar mer information på InfoFinlands sida Grundläggande utbildning.
Rådgivningsnumret 0800 9 8009 betjänar på finska och vid behov även på engelska eller svenska.
Familjemedlemmar till nordiska medborgare
Vid vissa universitet har olika examen olika namn.
Arbetarinstitutetfinska _ svenska _ engelska
Stödföreningen för unga invandrare R3 (R3 Maahanmuuttajanuorten tuki ry) hjälper ungdomar i frågor som rör utbildning och sysselsättning.
Dessutom kan du lista din arbetserfarenhet och utbildning i kronologisk ordning.
Du behöver inte ansöka separat om stödet, utan FPA betalar ut Vandatillägget (Vantaa-lisä) med hemvårdsstödet.
I vissa kommuner kan anmälan göras även på internet.
Barns och ungas problem
stöd för studerande
Om du vill kan du även be en stödperson att följa med.
Det öppna universitetet och de öppna yrkeshögskolorna har ett brett utbud av kurser också på engelska.
Information om presidentvalfinska _ svenska _ engelska
Karlebynejdens institutfinska _ svenska
Hjälp för invandrarmänfinska _ engelska
I Rovaniemi finns två hälsostationer:
FPA avgör om du har rätt att utnyttja socialskyddsförmånerna på basis av din ansökan.
studentexamen på finska eller svenska med ett godkänt vitsord i finska eller svenska som modersmål eller som andra språk
inledande kartläggning
I Finland finns en namnlag. Enligt den ska alla som har en hemort i Finland ha ett efternamn och 1–4 förnamn.
Navigatorn
Jämställdhetslagen förbjuder diskriminering på grund av kön.
Du kan studera vid flera olika läroanstalter: öppna universitetet (avoin yliopisto) eller öppna yrkeshögskolan (avoin ammattikorkeakoulu), sommaruniversitetet (kesäyliopisto), senioruniversitetet (ikäihmisten yliopisto), medborgarinstitut (kansalaisopisto), arbetarinstitut (työväenopisto) och folkhögskolor (kansanopisto).
Det är viktigt att känna till kollektivavtalet, eftersom det i Finland inte finns till exempel en lag om minimilöner, utan minimilönerna fastställs alltid enligt kollektivavtalet.
Klubbar för barnfinska _ svenska _ engelska
Ullavavägen 701, 68370 Ullava
Du hittar mer information om juridisk hjälp på InfoFinlands sida Behöver du en jurist?
innefatta internationell rörlighet i ett EU-program eller ett mångformigt program eller
I vissa undantagsfall kan man dessutom få medborgarskap på grundval av att man är född i Finland.
De hjälper både ungdomarna och föräldrarna i hedersrelaterade konflikter.
handledning och rådgivning för invandrare
Telefonnumret till jourmottagningen är 116 117.
Anmäl flyttningen till myndigheterna
Av plastförpackningarna tillverkas nya plastprodukter.
Att följa villkoren i hyresavtalet.
De flesta stöd ansöker man om av Fpa.
Din arbetsgivare behöver kortet för utbetalning av lön och för beskattningen.
Läs mer: Hobbyer för barn och unga.
Det betyder att till exempel sociala förmåner och lön minskar arbetsmarknadsstödets belopp.
Företagsfinland erbjuder en gratis telefontjänst där du får sakkunnig rådgivning om ditt företag har ekonomiska svårigheter.
Information om filmer och filmvisningarfinska _ svenska _ engelska
Du kan också kontakta A-kliniken.
Du kan även fråga om råd på rådgivningstjänsterna för invandrare.
År 1748 inleddes bygget av Sveaborgs sjöfästning på öarna utanför Helsingfors. (På finska Suomenlinna, "Finlands slott").
Ingen får särbehandlas till exempel på grund av kön, ålder, religion eller handikapp.
Barn i äktenskapet
Det finns även bidrag som du inte kan få om du inte bor stadigvarande i Finland eller har gjort det tidigare.
Du ska i allmänhet också betala de obligatoriska försäkringspremierna till Finland.
Service på svenska 0295 025 510
Lapplands universitet och Rovaniemi Steinerskola som är en privatskola.
Löneuppgifterna kan endast i undantagsfall anmälas med ett pappersformulär.
Om inget annat har avtalats i ditt hyresavtal räknas uppsägningstiden enligt lag från slutet av den månad under vilken du säger upp hyresavtalet.
Om du vill kan du även föda barnet på något annat sjukhus inom Helsingfors och Nylands sjukvårdsdistrikt (HNS).
Att uppgöra ett arbetsavtalfinska _ svenska _ engelska
Läs mer: Officiellt intyg om språkkunskaper.
Du kan ändå inte tacka nej till ett jobb som erbjuds till dig på grund av en utlandsresa.
Serviceboende ordnas för sådana handikappade personer som på grund av sitt handikapp eller sin sjukdom behöver hjälp för att klara av dagliga sysslor.
Flygtrafiken
i ett religiöst samfund som har rätt att förrätta vigsel
mån–tors kl. 8–16
Mer information om barns rättigheter i Finland hittar du på InfoFinlands sida Barn.
Om du är yngre än 30 år, kan du söka bostad hos Förbundet för ungdomsbostäder (Nuorisoasuntoliitto) och stiftelsen Nuorisosäätiö (Nuorisosäätiö).
Kostnader för ägarbostad
Hur påverkar det mitt uppehållstillstånd?
Din uppehållsrätt kan registreras om du studerar vid en läroanstalt som är godkänd i Finland.
Drygt en procent av befolkningen hör till den ortodoxa kyrkan.
Stöd för närståendevårdfinska _ svenska
Förutsättningen är inte att du är en infödd finsk medborgare, utan du kan också ha fått det finska medborgarskapet på ansökan.
I hälsorådgivningen beaktas hela familjen och ges särskilt stöd till den tidiga växelverkan.
Mer information om bostadsbidrag för pensionstagare hittar du på FPA:s webbplats.
Verksamhet för barnfamiljerfinska _ svenska _ engelska
Huvudregeln är att arbetsavtalet gäller tillsvidare.
Om du ansöker om dagvårdplats för första gången ska du använda den elektroniska ansökan.
Slott
Du kan också vända dig till Huvudstadens Skyddshem (Pääkaupungin Turvakoti).
De viktigaste besluten fattas på föreningsmöten som är öppna för alla medlemmar.
På familjerådgivningen kartläggs barnets situation så att barnet får den hjälp som det behöver.
Du hittar mer information om slotten och de guidade rundvandringarna på Museiverkets webbplats.
På familjeträningen får du också information om hur förlossningen sätter i gång och när det är dags att åka till sjukhuset.
Förlossningsavdelningen är öppen dygnet runt.
Flyktingen är i behov av internationellt skydd.
Hindersprövningen är obligatorisk och utan den kan vigseln inte förrättas.
Finlands riksdag beslutar hur många flyktingar som tas till landet.
De som har utexaminerats från en högskola eller ett universitet arbetar i många slags arbetsuppgifter.
På vintern är det kallt och snöar i Finland.
Läs mer: Graviditet och förlossning och När ett barn föds i Finland.
Medborgare i andra länder måste anmäla sig personligen vid TE-byrån.
Centria yrkeshögskolafinska _ svenska _ engelska
Den som har blivit förföljd på grund av sin sexuella läggning eller könsidentitet någon annanstans kan söka asyl i Finland.
linkkiFinlands Näringsliv EK:
Hemkommun i Finland
Det innebär att grundinformation om dig förs in i befolkningsdatasystemet.
Du kan även fylla i anmälan i magistraten.
Vem är barnets vårdnadshavare?
Mer information om barn vid skilsmässa finns på InfoFinlands sida Barn vid skilsmässa.
09 2313 9325 (mån.–fre. ll. 10–12)
Om du inte vill sköta bokföringen själv, kan du anlita en revisionsbyrå som sköter företagets bokföring åt dig.
Ingen skatt tas ut på barnbidrag.
Den inledande kartläggningen (alkukartoitus) hjälper dig att hitta lämpliga tjänster i din hemstad.
Även Karleby evangelisk-lutherska församlingssammanslutnings specialdiakoner erbjuder samtalshjälp vid missbruksproblem.
För arbetet under helgerna betalas högre lön.
Arbetsgivaren ingår vanligen ett skriftligt arbetsavtal med en ny anställd.
Omskärelse (ympärileikkaus) är alltid ett oåterkalleligt ingrepp.
linkkiFinlands Studentkårers Förbund:
en släkting som är bosatt i Finland har plötsligt insjuknat svårt eller avlidit,
Om du vill arbeta som företagare i Finland behöver du ett uppehållstillstånd för företagare.
Hälsostationerna har öppet vardagar kl. 8.00–16.00.
Boka en tid per telefon på numret (09) 4135 0501.
Grupperna i specialundervisningen är mindre än vanliga klasser.
A-klinikerna (A-klinikka) är vårdenheter där personer med missbruks- och beroendeproblem och deras närstående får stöd och hjälp. På A-klinikstiftelsens webbplats hittar du kontaktuppgifterna till A-kliniker runtom i Finland.
Väestöliitto erbjuder rådgivning och terapi för par på finska och engelska.
på finska 0295 020 500
Helsingfors rättshjälpsbyrå
Invånarna kan påverka stadens beslutsfattande redan då beslut bereds.
Hjälptelefon 0800 05058, mån.–fre. klockan 9–16
Nödsituationfinska _ svenska _ engelska
Du kan förlora din rätt till arbetslöshetsdagpenning för en viss tid om du själv har förorsakat arbetslösheten.
du är asylsökande och handläggningen av din ansökan är oavslutad
Då måste du i din ansökan be om att din information registreras i Finlands befolkningsdatasystem.
om du måste köpa receptbelagda läkemedel på apoteket för över tre månaders tid.
Detta betyder att man i situationen beaktar vad som är rimligt.
Läs mer: Barn vid skilsmässa.
Fundera också på vilka som är dina konkurrenter och hurdana produkter och verksamhetssätt de har.
Om flaggdagarna hittar du mer information på webbplatsen för Helsingfors universitets almanacksbyrå.
Innan du ansöker om utkomststöd ska du ansöka om de andra bidragen som du har rätt till (till exempel arbetslöshetsförsäkring, bostadsbidrag, pension, studiestöd, föräldradagpenning, sjukdagpenning, hemvårdsstöd eller underhållsstöd).
Service på finska 0295 025 500
Läroplikten är lagstadgad.
stödboende
Vid många yrkeshögskolor finns engelskspråkiga utbildningsprogram.
Ett samboförhållande kan utgöra ett hinder för att få uppehållstillstånd.
Vädret är svalt och ofta regnar och blåser det också.
har barnet rätt till familjepension om fadern dör.
Hälsostationerna har vanligen öppet från måndag till fredag kl. 310 1671.
På familjerådgivningen kan du diskutera familjens situation med de anställda.
Du ska alltid utreda din egen situation individuellt.
Barnbidrag betalas ut fram till dess att barnet fyller 17 år.
I EU-länderna finns några webbapotek där man kan lagligt köpa egenvårdsläkemedel.
Gemensam ansökan ordnas två gånger per år, på hösten och på våren.
Den vanligaste formen av människohandel är att tvinga någon till arbete utan lön eller under annars dåliga förhållanden.
Du får ett betyg för VALMA-utbildningen.
Vad ska jag göra?
Du kan boka en läkartid på din egen hälsostation.
Om alla uppgifter är korrekta, och det inte saknas några uppgifter, behöver du inte göra någonting.
koppleri.
Tfn (09) 816 42439
På Helsingfors stads webbplats hittar du information om skogen i Helsingfors och i närheten av Helsingfors.
Kontaktuppgifterna hittar du på organisationens webbplats.
Om du har elektriska värmeelement eller värmeaggregat hemma, lägg inte tyger, kläder eller något annat på dem.
Hälsovårdaren är på plats i skolan vissa dagar i veckan.
Korundifinska _ engelska
Staden ordnar boendetjänster till exempel för åldringar och handikappade, som har svårt att klara av de dagliga sysslorna utan hjälp.
När du kontaktar hälsostationen (terveysasema), bedömer en sjukskötare först din situation.
Man vet inte i förväg när förlossningen börjar.
Om du vill stanna kvar i Finland och registrera dig som invånare, ska du ha ett jobb eller ett aktivt företag, en studieplats, ett långvarigt familjeband eller tillräckliga medel.
Andra uppehållstillstånd för förvärvsarbete
Du kan även röra dig i naturen i Petikkos rekreationsområde.
Till en början var största delen av invånarna svenskspråkiga.
Kandidatstudierna pågår ungefär tre år, magisterstudierna ungefär två år.
Läs mer om kortvarigt boende på InfoFinlands sida Tillfälligt boende.
På InfoFinlands sida Studerande finns mer information för studerande som flyttar till Finland.
Mer information om skolorna i Vanda hittar du på Vanda stads (Vantaan kaupunki) webbplats.
Rådgivning erbjuds vid till exempel:
Information om möjligheter till fritidsaktiviteter hittar du på InfoFinlands sida Fritid.
Tfn 0295 016 620
Om du vill ha mer information om tjänster för äldre kan du kontakta seniorrådgivningen (seniorineuvonta).
Läs mer: Skilsmässa
Arbetsgivarna och arbetstagarna finansierar pensionsskyddet tillsammans.
Om man har hoppat av grundskolan, kan man avlägga grundskolans lärokurs också vid Eira vuxengymnasium (Eiran aikuislukio).
Ofta kan du skicka in ansökan och CV via arbetsgivarens webbplats.
De kan även köpa förskoleundervisningen till exempel av ett privat daghem.
Också sökandens inkomster beaktas, eftersom bostäderna främst är avsedda för personer med låga inkomster.
Det är fråga om barnkapning när
Du kan grunda ett företag i Finland oavsett ditt medborgarskap.
Med nationalpark avses ett över 1 000 hektar stort naturskyddsområde.
som inte står under förmyndarskap.
Grankulla stad har en egen begravningsplats i Kasabergsområdet.
Om du inte är medborgare i ett EU-land eller EES-land och inte heller familjemedlem till en medborgare i ett sådant land och du kommer till Finland för att studera i augusti 2017 eller senare, måste du betala terminsavgift för studierna.
Din hemkommun betalar assistentens lön.
Om du känner att du behöver hjälp omedelbart kan du kontakta den närmaste jourhavande hälsovårdscentralen eller sjukhusjouren.
Anmälan till grundskolan ska göras på förhand.
Mer information om högskolorna i Esbo och Helsingfors hittar du på städernas webbplatser.
Skilsmässoansökan(pdf, 100 kb)finska _ svenska
Finland som flykting utarbetas en inledande kartläggning och integrationsplan för dig vid utlänningsbyrån.
På sommaren är nätterna för ljusa för att man ska kunna se norrsken.
När du ansöker om tillstånd tas dina fingeravtryck för det biometriska uppehållstillståndskortet.
Den utländska partnern behöver dessutom ett identitetsbevis, ett civilståndsintyg (ogift, skild, änka/änkling) och ett Apostilleintyg för dessa.
I brådskande nödsituationer ska du ringa nödnumret 112.
Sändaren ska inhämta ett skriftligt tillstånd för offentlig visning av videoklippet av samtliga personer som uppträder i videoklippet och kan identifieras, samt av de personer som medverkat i framställningen av videoklippet.
Information och råd om var du kan få hjälp med olika slags problem i arbetslivet hittar du på InfoFinlands sida Problem i arbetslivet.
Utländskt körkort i Finlandfinska _ svenska _ engelska
Läs mer om förutsättningarna på sidan EU-medborgare.
verksamhetslokaler
Specialpedagogik i förskolanfinska _ svenska
Karlebynejdens institut erbjuder barn och unga olika former av hobbyverksamhet, exempelvis i konstämnen och musik.
Automaten skriver ut en parkeringsbiljett som du placerar innanför bilens vindruta så att hela parkeringsbiljetten kan läsas från utsidan.
Språkcentret vid Lapplands universitet ordnar kurser i finska språket på engelska.
linkkiTeaterinfo Finland:
I Vanda finns flera yrkes- och amatörteatrar.
Om bostaden är byggd med statsstöd, kan du ansöka om
Folkhögskolornas ansökningspraxis och ansökningstider varierar.
Alla arbetstagare ska behandlas jämlikt och lika.
Var aktiv.
disponera över sin egendom
Barnets för- eller efternamn kan inte bytas utan barnets tillstånd.
Teckna en tillräckligt omfattande sjukförsäkring i ditt hemland
När du går till magistraten ska du ta med dig
Den offentliga tandvården
Du får förvärvsarbeta i Finland om det har gått tre månader sedan du lämnade in din asylansökan och du har ett giltigt pass eller någon annan resehandling som du har företett till myndigheten när du sökte asyl.
I Finland bestäms arbetstagarnas rättigheter enligt arbetslagstiftningen och kollektivavtalen (työehtosopimukset).
Införsel av flyttsaker till Finlandfinska _ svenska _ engelska _ ryska
linkkiSHVS:
Farsdag firas i Finland den andra söndagen i november.
Att köra bil och parkera
Spara arbetsintyg för eventuella granskningar.
Om du behöver en tillfällig barnskötare hem, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Mer information hittar du på webbplatsen.
De är alltså avsedda för alla invånare i staden.
Det är bra att fundera på vilket språk du vill registrera för ditt barn.
Försök att enas om saken med hyresvärden innan avtalet hävs.
Information om utkomstskyddet för arbetslösafinska _ svenska _ engelska
Grundläggande utbildning
Hyresbostäder i Rovaniemifinska
Makar har giftorätt till varandras egendom.
Sjukdagpenningfinska _ svenska _ engelska
Du kan delta i tävlingen fram till den 1 december 2013.
Ofta är ansökningstiden fortlöpande.
Information om utsökningfinska _ svenska _ engelska
Ounasrinteentie 22
Sjöstöveln 1 A
NewCo Helsinki erbjuder rådgivning och hjälp med att starta eget företag på finska, svenska, engelska, ryska, arabiska, estniska, tyska och italienska.
Hälsocentralsjourenfinska _ svenska _ engelska
Även klädskåp och skåp i hallen ingår vanligtvis.
Tjänsterna inom kommunernas ungdomsarbete är avsedda för barn och unga vuxna.
Garantipensionen betalas inte om du flyttar utomlands för över ett år.
Det behövs minst tre personer för att grunda ett andelslag.
I Helsingfors finns Global Clinic, där personer som vistas i Finland utan tillstånd kan få primärhälsovård.
För hormonella preventivmedel behöver du ett läkarrecept, som du får till exempel från hälsostationen eller av en privat gynekolog.
Att meddela hyresvärden om du upptäcker sådana fel i bostaden som hyresvärden ansvarar för.
Om du har bevis på hot och trakasserier är det bra att spara dem.
Den förälder som inte bor med barnet betalar underhållsbidrag till den förälder hos vilken barnet bor officiellt.
Finska som andra språk i den grundläggande undervisningenfinska
Du hittar information om den finländska kulturen på InfoFinlands sidor Finländska seder och Den finländska arbetskulturen.
Förbered dig på företagande
I ditt bostadsområde arbetar dessutom stadens kontaktperson, stadslotsen (stadiluotsi), som kan hjälpa dig att föra vidare ditt förslag.
moderns efternamn eller
De som arbetar med barnen är utbildade pedagoger inom småbarnsfostran och barnskötare.
Om du har frågor om den grundläggande utbildningen kan du även kontakta stadens undervisningstjänster.
Du kan endast använda faderskapspenningdagar för vård av ett barn under två år.
Vårdnaden är inte beroende av vem barnet bor med.
I nästan alla högskolor erbjuds dock även undervisning på engelska.
Finlands första universitet
linkkiFörbundet för ungdomsbostäder rf: Boendehandbok för ungdomarfinska
Bland annat vid månadsskift och på veckoslut är flyttfirmorna alltid upptagna.
uppehållstillstånd som är giltigt i minst ett år; eller
Stöd vid ekonomiska problem
Annan viktig information om boendet i Finland finns på InfoFinlands sida Boende.
Även om du klarar dig i många dagliga situationer på engelska kräver de flesta arbetsgivare att du kan finska eller svenska.
Arbetsavtalet för en gravid kvinna får inte hävas och hon får inte diskrimineras på grund av sin graviditet.
Religiösa samfundfinska _ svenska _ engelska
Utredning över samboskap (om du är sambo med EU-medborgaren och ni inte har gemensam vårdnad om barn)
Handikappbidragets storlek beror på hur svårt ditt handikapp är.
Fråga mer om distansstudier vid ditt eget gymnasium.
Du kan ersätta statsförvaltningens språkexamen med vissa andra studier.
Tredjelandsmedborgare äe medborgare i annat land än de nordiska länderna, EU-länderna, Liechtenstein eller Schweiz.
registrerat dig som arbetslös arbetssökande vid arbets- och näringsbyrån
Tfn 040 559 6564
Erkännande av faderskap
Invandrare får hjälp med jobbsökningen vid Lapplands arbets- och näringsbyrå (TE-byrån).
rätt att rösta i presidentval, riksdagsval och folkomröstningar då man fyllt 18 år.
Tfn 010 235 1450 (kundtjänst)
Var noga när du fyller i ansökan.
Tilläggsövningar till läroboken Hyvin meneefinska
Du kan inte söka till en yrkesinriktad vuxenutbildning i den gemensamma ansökan.
Om ni inte kan komma överens om hur ni ska dela upp egendomen, kan vem som helst av makarna kräva egendomsfördelning, det vill säga bodelning (ositus).
Där kan eleverna höja sina vitsord och fundera på vilket studieområde de är intresserade av.
Begär tillståndet skriftligt.
För gymnasium förberedande undervisningfinska _ engelska
ditt pass där ditt uppehållstillstånd syns
Jämställdhetslagen förbjuder diskriminering på grund av kön.
Läs mer: Problem i äktenskap och parförhållande
Öppet
små plastleksaker och bruksföremål i plast såsom disk- och tandborstar.
Vuxengymnasiet är i huvudsak avsett för personer som har fyllt 18 år.
Mångkulturell barndagvård
Kommunerna ordnar medicinsk rehabilitering till exempel vid hälsovårdscentraler och i sjukhus.
Hindersprövningen görs i magistraten (maistraatti).
Fpa om du flyttar utomlands permanent eller vistas utomlands mer än tre månader.
Arbete som freelancer innebär att du arbetar för flera uppdragsgivare utan fast anställning.
Kontrollera på institutets webbplats vilka kurser som är aktuella.
Därefter larmar han eller hon hjälp.
Studierna är avgiftsbelagda.
Lokaltrafiken trafikeras vanligtvis med bussar.
linkkiArbets- och näringsministeriet :
Varje barn har rätt till en god och trygg barndom.
Om misstanken är befogad, kan det beslutas att umgänget ska ske under socialmyndigheters uppsikt.
Volontärarbeteengelska
Inom den grundläggande utbildningen (ungdomar och vuxenstuderande)
Om det finns minst tre elever som befriats från religionsundervisningen och deras föräldrar kräver detta, ordnas undervisning i elevernas egen religion.
Sjukvård för utlänningar i Finlandfinska _ svenska _ engelska
avläggande av delar av ovan nämnda examina.
Boendevardag
Luckan Integration är en rådgivningstjänst, som erbjuder personlig rådgivning för invandrare och anordnar bland annat evenemang och grupper relaterade till jobbsökning.
Mattsgatan 7
Ofta kan du få betalningstiden förlängd.
Om du ska flytta till Finland för studier måste du ta hand om följande:
Socialrådgivningfinska _ svenska
Ungdomarna har många möjligheter att påverka.
Fasta hjälpmedel kan till exempel vara olika typer av lyftanordningar samt brandvarnare och dörrklocka för hörselskadade, där ljudet har ersatts med lampor.
Kontaktuppgifterna till barnatillsyningsmannen hittar du på Vanda stads webbplats.
Till exempel ger ett uppehållstillstånd på grund av familjeband mer omfattande rätt att arbeta än ett tillstånd som beviljats på grund av studier.
Fullmäktige väljs vart fjärde år genom kommunalval.
Du kan också komma utan tidsbokning för att prata om din situation, måndag till fredag kl. 9–11 och onsdagar kl. 16–20.
De flesta lagarna från den svenska tiden fortsatte att gälla.
Beslutsfattandefinska _ svenska _ engelska
Det är dock många som ansöker om stadens bostäder och endast en liten del av de sökande får en bostad.
Du kan idka båda grenarna på egen hand när du väl lärt dig grunderna.
Arbete ger dig åtminstone delvis rätt till den sociala tryggheten i Finland
skuldrådgivning
Detta är dock inte alltid möjligt.
Den tillfälliga barnpassningshjälpen är avgiftsbelagd.
Vanligen ger man inte varandra presenter på arbetsplatserna.
Du kan ansöka om lånegaranti vid Takuusäätiö om du behöver ett banklån för att betala dina skulder.
_ danska
du är arbetslös arbetssökande eller
ett barn under 16 år som är bosatt i Finland förs utomlands utan vårdnadshavarens tillstånd
Många finländare badar bastu varje vecka.
Om du upptäcker att du själv eller en närstående får allt svårare att komma ihåg saker, kan du kontakta hälsostationen i ditt område och boka en tid hos läkaren.
Läs mer: Problem i äktenskap och parförhållande.
När du är gravid kan FPA betala ut moderskapspenning (äitiysraha) till dig.
Lapplands universitet och Rovaniemi Steinerskola som är en privatskola.
Läs mer om tolktjänsterna på InfoFinlands sida Behöver du en tolk?
Till vissa utbildningsprogram antas endast en liten del av sökandena.
De ordnar verksamhet under 2–5 dagar i veckan med tyngdpunkt på fredagar och lördagar.
Beskattningsbeslut
Polisen anmäler brott som begåtts av barn under 18 år till föräldrarna och barnskyddsmyndigheten.
Ungdomsgården Vinge
Du måste även låta översätta handlingarna till finska, svenska eller engelska om de är på något annat språk.
Företagare måste ändå ordna företagshälsovård för sina anställda.
Fakturan kan uppgå till flera tiotusentals euro.
Du kan även boka tid hos en privat gynekolog.
Om det inte är möjligt fattar läkaren beslut om kejsarsnitt.
Att åka skidor är en av de populäraste vintersporterna i Finland.
Du kan anmäla dig via Internet om du har finländska webbankkoder.
Kontaktuppgifter:
Om den unga begår ett brott kan han eller hon åtalas och dömas för det.
När du öppnar ett bankkonto behöver du ett pass eller någon annan officiell identitetshandling.
Information om hobbyverksamheter för barn och unga finns på stadens webbplats.
Läget som granne till huvudstaden Helsingfors har varit viktigt för Vanda.
Ansökan till förskoleundervisningfinska _ engelska
Barnet kan vid behov även få ett skolgångsbiträde (koulunkäyntiavustaja).
Ansökan om moderskapsunderstöd och moderskapspenning
EU-länderna, EES-länderna och Schweiz
Hjälp med ekonomiska problemfinska _ svenska _ engelska
Också nya elever har rätt till denna stödundervisning.
Bussar
Kontaktuppgifter till FPAfinska _ svenska _ engelska
Därtill finns det intervjuer, diskussioner och skriftliga uppgifter.
På en finländsk arbetsplats övervakar chefen inte de anställdas arbete hela tiden.
Läs mer: Andra studiemöjligheter.
Läs mer om LUVA-utbildningen på InfoFinlands sida Förberedande gymnasieutbildning.
Elever som har finska som modersmål lär sig svenska i skolan.
Se till att din bostad hålls i gott skick.
Läs mer på InfoFinlands sida Den sociala tryggheten i Finland.
Haartmanska sjukhuset
Den som säljer en bostadsaktie är vanligen ansvarig för fel under två år.
När ett barn föds till familjen kan modern eller fadern enligt lag stanna hemma för att ta hand om barnet.
I första hand försöker man använda öppenvården alltså att barnet bor tillsammans med sin familj.
hushållsavdrag
Giltigt pass
Be om tips till jobbsökningen och hjälp med att skriva ansökningar av andra.
Med underuthyrning avses att hyresgästen hyr ut en del av bostaden till en annan person.
Telefon: 029 566 1270
ett intyg på vederlagets belopp och bostadslånet (ägarbostad)
På den internationella träffpunkten Trapesa kan du delta i en samtals- och inlärningsgrupp på finska.
Lapplands läroavtalscenter
Åbovägen 150
68370 Ullava
Staden har åtagit sig att sörja för integritetsskyddet för användarna av stadens webbtjänster.
Samarbetsprojektet Versofinska
Finska ortodoxa kyrkanfinska _ svenska _ ryska
Ofta kan du även skicka in en öppen ansökan via företagets webbplats.
Om du råkar ut för problematiska situationer på arbetsplatsen ska du först kontakta din chef.
vistas i Finland av någon annan orsak än studier.
Begravningsbyråerna säljer också kistor och sköter enligt avtal och de anhörigas önskemål även allt annat som rör begravningen.
En engelskspråkig förteckning över konventionsstaterna finns på webbplatsen för internationella domstolen i Haag.
Adress: Brunnsgatan 1 (Helsingfors huvudjärnvägsstation)
jobbsökningsförmåga och planerar sin framtid.
Arbets- och näringsbyråerna tillhandahåller till exempel följande tjänster:
Kontaktuppgifter och tjänsterfinska _ svenska
Du kan till exempel få hjälp med psykiska problem och missbruksproblem samt hjälp att sluta spela.
Kontakta Karleby stads förskoleundervisning för information om specialsmåbarnspedagogiken.
Om du på grund av ditt handikapp behöver till exempel en speciell dator eller särskilda hushållsapparater kan du få understöd för detta vid socialbyrån i din hemkommun.
Köpcentret Grani
Asylsökanden kan beviljas flyktingstatus om han eller hon har befogade skäl att frukta förföljelse i sitt hemland på grund av ras, religion, nationalitet, tillhörighet till en viss samhällsgrupp eller på grund av sin politiska uppfattning och då sökanden på grund av detta inte kan återvända till sitt hemland.
Om du är sjukförsäkrad i Finland, får du ett FPA-kort.
Ensamkommande barn(pdf, 674)finska _ svenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ persiska _ arabiska _ kurdiska
Ofta kan du även fylla i och skicka blanketten på kommunens webbsida.
_ slovakiska
öppettider:
I Finland ska barnen delta i förskoleundervisning under ett års tid innan läroplikten börjar.
Utan dem är det mycket svårt att ta sig upp ur en vak.
I nödsituationer får du vård även om du inte har en hemkommun i Finland.
Hälso- och sjukvårdstjänster lämnas på finska och svenska i Finland.
Hos dessa organisationer kan du få råd och hjälp till exempel vid ansökan om tjänster.
I biblioteket kan du också använda dator.
Att anmäla sig som kund
Information om utbytesprogrammetengelska
Magistraten undersöker om det finns hinder mot äktenskapet utifrån de uppgifter som finns registrerade i Finlands befolkningsdatasystem.
Det förutsätter att modern eller fadern varit anställd hos samma arbetsgivare minst sex månader under det senaste året.
Man söker till yrkesutbildning i den gemensamma ansökan.
NEJ: farligt avfall
Ansökningen kan tas för behandling först när du besökt beskickningen eller tjänstestället.
Vistelse i skyddshemmet är kostnadsfritt.
Rådgivningen på olika språk:
Om föräldrarna inte är gifta kan barnet få antingen moderns eller faderns efternamn, om faderskapet har fastställts.
I Finland finns åtta kommunala tolkcentraler (tulkkikeskus).
På Vanda konstmuseum ordnas växlande utställningar med inhemsk och utländsk modern konst.
vikariat
Magistraten i Västra Finland
Du kan avlägga utbytesstudier via olika program.
Asylsökande som inte beviljas flyktingstatus kan ändå få uppehållstillstånd i Finland på någon annan grund.
Om du vet att du kommer att bli sen till arbetet ska du tala om det för din chef.
Om du på grund av ditt handikapp inte kan använda kollektivtrafiken kan du ha rätt till färdtjänst (kuljetuspalvelu).
Till arbets- och näringsbyråns (työ- ja elinkeinotoimisto) kurser i finska eller svenska ansöker du via arbets- och näringsbyrån.
Läs mer om prövning av äktenskapshinder på InfoFinlands sida Prövning av hinder mot äktenskap.
Att se till att hyresbostaden hålls i ett gott skick.
Yrkesutbildning
På InfoFinlands sida Utkomstskydd för arbetslösa får du mer information om vem som har rätt till utkomstskydd för arbetslösa.
Högskolor som erbjuder SIMHE-tjänsterfinska _ engelska
Till exempel ändrade familjeförhållanden eller att du börjar arbeta kan påverka din rätt till FPA:s förmåner.
har förvärvat sitt medborgarskap på grund av faderns finska medborgarskap och faderskapet upphävs.
Grunderna för antagning av studeranden beror på utbildningen.
På så sätt kan man bevisa att lönen verkligen har betalats till dig.
Ofta krävs det även att personen bosatt i Finland ska ha tillräckliga medel för att försörja en familjemedlem som flyttar till Finland.
Det finns inga egentliga nationella prov.
Du kan också vända dig till rådgivningstjänsten för invandrare i din kommun.
Glas (lasi)
ägna dig åt båtliv, simma och tvätta dig i sjöar och vattendrag samt färdas på isen.
Filmerfinska _ svenska _ engelska
På rådgivningsbyrån följer en hälsovårdare ditt hälsotillstånd och babyns hälsa.
Via beskickningen kan du ofta uträtta till exempel följande ärenden:
kan på ett pålitligt sätt styrka sin identitet
Blandavfall (sekajäte) eller övrigt avfall
Du kan studera vid en öppen yrkeshögskola även om du inte har någon examen.
För att barnet ska kunna få uppehållstillstånd måste hans/hennes uppehälle i Finland vara tryggat, till exempel genom förälderns löneinkomster.
Skatteförvaltningen
Äktenskapet är alltid ett frivilligt val som ingen kan tvingas till.
Semester, studier eller arbete under arbetslösheten
Kontaktuppgifter:
Referenser – Du kan lägga till namnen på personer som har lovat att rekommendera dig för arbetsuppgiften.
Frågor som rör skolgången för ett handikappat barn kan du ställa till skolväsendet (opetustoimi) samt till servicehandledaren för skolelever (koululaisten palveluohjaaja).
Båda pensionerna kan sökas hos Fpa.
Vanligast är att äktenskapsförordet fastställer att ingendera maken har rätt till den andras egendom.
Bibliotek och öppettiderfinska _ svenska _ engelska _ ryska
Yrkesutövarnas och företagarnas arbetslöshetskassafinska _ svenska _ engelska _ ryska _ estniska
Invandrarrådgivarna i din kommun i Finland
Till exempel studerande har denna möjlighet.
Om du vill ha en religiös vigsel kommer du överens om detta med ett religiöst samfund.
Studier som hobby, Arbetskraftsutbildning
På din lön eller annan inkomst har det innehållits skatt utgående från skattekortet.
arbetsförsök
Varje sökandes livssituation behandlas individuellt när FPA fattar beslut om bidrag.
När du funderar på om det är finska eller svenska som du borde lära dig ska du beakta vilket språk som talas på din hemort och i din näromgivning.
Du kan använda svenska med statliga myndigheter, till exempel FPA eller TE-byrån.
Gymnasiestudierna pågår vanligen tre år.
växtodling
Skattebyrån
Om du inte kan komma överens om löneutbetalningen med din arbetsgivare måste ärendet avgöras i domstol.
Tfn 029 5645 000
Du kan registrera dig som arbetslös arbetssökande elektroniskt
Också asylsökande kan använda tjänsterna vid mödrarådgivningen.
Hurdana ljud är tillåtna i ett höghus?
Läs mer: Registrering som invånare.
Alla kan själv välja var de vill bo och fritt röra sig i Finland.
Bussar
Mer information finns på InfoFinlands sida Översättningar
Remiss för hemsjukvården skrivs av läkare.
linkkiFFC:
Diskutera först med din läkare inom företagshälsovården och din arbetsgivare om möjligheten att söka partiell sjukdagpenning.
Kivenkolo
Lekparkerna och familjehusen ordnar vården av barnen under den tid kursen varar.
I Finland ordnas också många teaterfestivaler.
Legaliserade födelseattester för dina barn i original (om du har barn under 18 år som flyttar till Finland)
Könsstympning av flickor är ett brott i Finland.
Hjälp i frågor om utbildning
Du får rådgivning på finska och engelska.
Hyresgaranti
Ring fastighetsskötseln som ditt bostadsaktiebolag har avtal med.
Studierna vid öppna högskolor är inte heltidsstudier.
Du ska ändå lämna in din ansökan i den egna kommunen.
Heminkvartering
en ägarbostad
FPA ersätter högst 80 terapibesök om året och högst 200 besök under tre år.
Vanligtvis ska du sortera avfallet hemma innan du gör dig av med det.
Om båda föräldrarna arbetar, har barnet rätt till småbarnspedagogik på heltid.
Du kan begära hindersprövning på vilken magistrat som helst.
Du kan skicka uppgifterna om din affärsverksamhetsplan och erforderliga handlingar till Business Finland på elektronisk väg.
Säkerhetsbranschen
Av dem är cirka 2,8 procent svenskspråkiga och 11 procent har något annat modersmål än finska eller svenska.
När myndigheten har mottagit din asylansökan, hänvisas du till ett mottagningscenter.
Dessa bostäder hittar du på studentkårens webbplats.
Om intyget har utfärdats av en myndighet i ett EU-land och åtföljs av blankett EU 2016/1191, behöver intyget inte översättas.
Underhållsbidrag
Information om räntestödetfinska _ svenska _ engelska
Sökning av hyresbostäderfinska _ engelska
Skolhälsovårdenfinska _ svenska
Skatteförvaltningens riksomfattande telefontjänst: 029 497 050
Dessa arbetsgivare ger garanti om en arbetsplats.
Finländarna är också aktiva paddlare och seglare.
Sök till gymnasiet i den gemensamma ansökan till andra stadiet i februari-mars.
Lägg inte skräp, mat eller kemikaler i avloppet (WC:n).
Man kan också söka skilsmässa ensam.
Integrationsutbildning
Ta kontakt med din läkare, företagsläkare eller FPA.
Du kan lämna in din ansökan om identitetskort på vilken av polisens tillståndsenheter som helst.
Polisen ser till att dödsorsaken fastställs och anmäler dödsfallet till Befolkningsregistercentralen (Väestörekisterikeskus).
Kom ihåg att alltid begära ett intyg när du haft ett jobb, avlagt en praktik eller studerat.
Om du vill ansöka om finskt medborgarskap behöver du ett officiellt intyg över dina kunskaper i finska eller svenska.
Ryssland ockuperade Helsingfors två gånger på 1700-talet när Sverige och Ryssland var i krig.
Om den avlidne har arbetat eller varit företagare i Finland kan dennes efterlevande få familjepension från arbetspensionssystemet.
Du kan kontakta diskrimineringsombudsmannen byrå om du har råkat ut för diskriminering eller upplever att du har bemötts rasistiskt eller osakligt på grund av ditt etniska ursprung eller för att du är utlänning.
linkkiRovaniemi stads ungdomstjänster:
Läs mer: Våld
en uppskattning av dina inkomster för hela året
Naturobjekt i Esbofinska _ svenska _ engelska
Ring inte nödnumret om det inte är fråga om en nödsituation.
Legaliserat äktenskapsintyg i original (om du är gift)
Också sambor kan få hjälp med att komma överens om saker och ting, till exempel genom medling i familjefrågor.
tfn 016 322 4600
De behöver till exempel inte be om tillstånd av släktingar.
I Finland har alla möjlighet att få avgiftsfri företagsrådgivning.
Genom fristående examen kan du avlägga
Mer information om medborgarskapsansökan och om annat som rör medborgarskap får du på Migrationsverkets webbplats.
Elektroniskt responssystemfinska _ svenska _ engelska
Du får själv bestämma om du tar ut alla faderskapspenningdagar eller bara en del av dem.
Östanvindsvägen 1 A
folkpensionen, garantipensionen och andra bidrag för pensionärer
Dagvård fås på finska och på svenska.
På TE-byråns jobbsajt finns tusentals arbetsplatser runt om i Finland.
Du kan ansöka om Karlebystödet om den ena av föräldrarna vårdar samtliga av familjens barn under skolåldern i hemmet.
Du kan kontakta Brottsofferjouren per telefon eller via chatten eller besöka servicepunkten.
Observera att alla beskickningar inte erbjuder samma tjänster.
Vid magistraten kan du få en finsk personbeteckning, om du inte fick den redan i samband med att du beviljades uppehållstillstånd eller din uppehållsrätt för EU-medborgare registrerades vid Migrationsverket.
Kriscentret Monikas hjälptelefon är avsedd för invandrarkvinnor.
Trafiken
Läs mer på InfoFinlands sida Nordisk medborgare.
Dra dig alltså inte för situationer där du har möjlighet att tala finska eller svenska.
En utvecklingsstörning gör det svårare att lära sig och förstå nya saker.
Du kan åka till Böle eller beställa material till ditt eget närbibliotek.
På magistratens webbplats finns mer information om registreringen av utlänningar.
Införsel av läkemedel till Finlandfinska _ svenska _ engelska
Tandvården
Före äktenskapet ska ni tillsammans skriftligt begära hindersprövning (esteiden tutkiminen).
Offentliga hälsotjänster tillhandahålls vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Om du vistas i Finland mer än tre månader, behöver du ett registreringsintyg för EU-medborgare (Unionin kansalaisen rekisteröintitodistus).
Alla som bor i Finland måste följa Finlands lag.
I Vanda finns jourmottagningen på Pejas sjukhus (Peijaksen sairaala).
är minst 18 år gammal
Om ett sjukt barn behöver läkarhjälp eller uppsöka hälsovårdare ska du kontakta hälsostationen (terveysasema) eller en privat läkarstation i din hemkommun.
Säg inte upp din försäkring.
Den egendom som maken har vid ingående av äktenskap eller förvärvar under äktenskapet förblir hans tillhörighet.
Arbetsgivaren kan också ordna sjukvårdstjänster för sina anställda.
Finlands grundlagfinska _ svenska _ engelska _ ryska _ franska _ spanska _ tyska
Det finns emellertid många sökanden till stadens bostäder och bara en liten del av alla sökanden får en bostad.
Advokaterfinska _ svenska _ engelska
Notera att du måste besöka magistraten personligen.
Information om förmedling i familjefrågorfinska _ svenska _ engelska
Helsingfors historia
Vårdpenning betalas bara för ett barn i taget och är skattepliktig inkomst.
I Helsingfors finns SERI-stödcentret som är avsett för offer för sexuellt våld.
Familjeförmåner utomlandsfinska _ svenska _ engelska
Förvärvsinkomsten ska vara ungefär lika stor som företagarens genomsnittliga lön skulle vara om han eller hon skulle utföra liknande arbete som anställd.
Bearbeta – remixa, transformera, och bygga vidare på materialet för alla ändamål, även kommersiellt.
Till exempel kan föräldrar få föräldradagpenning endast om de har bott i Finland minst 180 dagar före barnets beräknade förlossningsdatum.
Om familjen inkomster är mycket låga, kan småbarnspedagogiken vara kostnadsfri för familjen.
Läs mer på InfoFinlands sida Företagshälsovård.
Kulturevenemangfinska _ svenska _ engelska
Du behöver inget uppehållstillstånd i Finland.
Personalen vid Navigatorn hjälper dig om du inte har något arbete eller en studieplats.
Registrerat parförhållande
Tfn: (09) 8392 4202
linkkiNorra Finlands tolktjänst:
Gym för äldrefinska
Ett recept som du skaffat utomlands är inte giltigt i Finland.
Ange en länk till webbplatsen InfoFinland.fi och nämn licensen CC BY 4.0.
linkkiArbets- och näringsbyråns tjänster:
I sista hand avgörs ärendet i tingsrätten.
Information om att öppna ett bankonto finns på InfoFinlands sida Vardagslivet i Finland.
Under VALMA-utbildningen får du kunskap och färdigheter som hjälper dig i dina senare yrkesinriktade studier.
Om du kommer till Finland från utlandet för att arbeta, behöver du en finsk personbeteckning.
Tolken är en neutral, utomstående person som varken är på din eller på myndighetens sida.
Giltigt pass
Arbete och studier
Läs mer om arbetsavtalet på InfoFinlands sidor Att komma överens om anställningsvillkoren och Innehållet i arbetsavtalet.
Fråga mer hos FPA:s center för internationella ärenden.
Rätten till barnbidrag upphör.
Observera att tjänstestället inte kan ge rådgivning om tillståndsärenden.
På många arbetsplatser har man flexibel arbetstid och man kan komma till arbetet till exempel mellan klockan 7 och 9 och gå hem mellan klockan 15 och 17.
linkkiSAMOK:
Läs mer: Problem i äktenskap eller parförhållande.
Det är inte möjligt att säga upp ett tidsbestämt avtal under dess giltighetstid.
Arbetsavtalslagen beskriver vilka orsaker som är godtagbara för uppsägning.
Intyget över hindersprövningen är i kraft fyra månader.
Förfrågningar om hyresbostäder på Rovaniemi stads område kan ställas direkt till fastighetsägare eller till bostadsförmedlingar.
Ytterligare information om yrkesutbildningfinska _ svenska _ engelska
Byråarbetare
Klimatet i Finland är kallare än i många andra länder.
Sexualhälsa
Barnen börjar i förskoleundervisningen vanligen vid sex års ålder och grundskolan vid sju års ålder.
Du blir också tvungen att betala ränta på kvarskatten efter en viss tid.
Domstolen kan även begära en utredning av kommunens socialväsen.
Teckna försäkringar
för att arbeta,
Ett samboförhållande upphör när parterna inte längre bor på samma adress.
Tfn (09) 8392 0071
Rådgivningsbyråerfinska _ svenska _ engelska
I Finland beskrivs språkkursernas nivåer på olika sätt.
Examen på utmärkt nivå kan endast avläggas i Helsingfors.
barn
Läs mer om beskattningen i Finland på InfoFinlands sida Beskattning.
Utöver den betalda semesterna kan du ansöka om obetald ledighet.
Om du har ekonomiska problem kan du be om råd hos Mellersta Österbottens social- och hälsovårdssamkommun Soites enheter för socialarbete eller utkomststöd, tfn 040 806 5095 eller tjänstestyrningen, tfn 040 806 5093.
Vid medborgarinstitutet kan man till exempel skapa konst, göra handarbeten, laga mat, dansa eller motionera.
studentexamen eller en motsvarande examen i ett annat land
Handikappade personer
När faderskapet har fastställts
InfoFinlands
Till exempel omfattar nivå A1 kurserna A1.1, A1.2 och A1.3 och nivå A2 kurserna A2.1 och A2.2.
Avfallshantering för bostaden finska _ svenska
Social- och krisjouren
Föräldrarna kan förvänta att flickor beter sig på ett annat sätt än pojkar.
På Helsingfors stads webbplats hittar du en lista över de daghem och skolor som ger förskoleundervisning.
Anvisningar för dig som ska grunda ett café eller en restaurang finska _ engelska
Serviceguide för seniorer(pdf, 1,8 MB)finska _ svenska
Om du inte är medlem i ett fackförbund, kontakta till exempel arbetarskyddsmyndigheterna.
Hälsostationen har öppet vardagar kl. 8.00–16.00.
Minderåriga asylsökande
Man kan insjukna i typ 2-diabetes (diabetes) i vilken ålder som helst men ofta insjuknar man i pensionsåldern.
Prepaid-abonnemang kan köpas till exempel i R-kiosker, en del snabbköp och på Internet.
Du kan kontrollera hos regionförvaltningsverken eller på Företagsfinlands webbplats om du behöver ett tillstånd för ditt företag.
Om du har fått för lite lön, ska du be din arbetsgivare att rätta till löneutbetalningen.
I hälso- och sjukvården av barn under skolåldern får man hjälp av rådgivningens hälsovårdare och läkare.
Ibland kan föräldrarna inte sörja för barnets välfärd.
sophämtning
Familjerågivningscentralen
Om du eller din familj inte har tillräckliga inkomster eller tillgångar för den nödvändiga dagliga försörjningen kan du söka grundläggande utkomststöd hos FPA.
Hjälpmedel för att röra sigfinska _ svenska
linkkiKulturhuset för barn och unga Fernissan:
Mer information hittar du på Asuntosäätiös webbplats.
Studentskrivningarna (ylioppilaskokeet) skrivs oftast i slutet av studierna.
Du kan flytta in i bostadsrättsbostaden när du har gjort bostadsrättskontraktet och betalat bostadsrättsavgiften.
Du kan skaffa könumret via internet.
En grundskolebaserad utbildning varar i cirka tre år.
Den närmaste flygplatsen är Helsingfors-Vanda flygplats.
Läs mer på InfoFinlands sida Medier i Finland.
Esbo stad betalar ett kommuntillägg till de familjer som vårdar ett under treårigt barn i hemmet.
hälsotillstånd
Hjälptelefon: (09) 276 62 899
På museet finns Renlunds samling av finländsk konst från guldåldern och tillfälliga utställningar i en kulturhistorisk miljö.
Teknik och kommunikation
Tfn (09) 4777 180 (24h)
Med energiavfall avses bl.a.:
En anställd vid arbets- och näringsbyrån (työ- ja elinkeinotoimisto) upprättar en inledande kartläggning (alkukartoitus) och en integrationsplan (kotoutumissuunnitelma) tillsammans med dig när du registrerar dig som arbetssökande.
Boka tid per telefon på nummer (09) 413 50 510.
Information om uppehållstillståndfinska _ svenska _ engelska
religion
Läs mer på InfoFinlands sida Förberedande gymnasieutbildning.
Du kan söka svenskspråkig yrkes- och gymnasieutbildning samt förberedande utbildning före dessa via tjänsten Opintopolku.fi.
Med statens lokalförvaltning avses de myndigheter som sköter statliga ärenden i en viss region.
Hyresvärden kräver att jag betalar hyra även för juli.
Fackförbundets medlemmar kan delta i utbildning och fritidsaktiviteter som förbundet ordnar.
Finländarna ser sig själva som västeuropéer, eftersom tiden som en del av det svenska riket knöt finländarna starkt till det västliga kulturarvet.
Många finländare åker gärna till stugan på midsommaren.
Sjukhusgatan 3 (Räckhals gård)
I vissa fall ersätter Kela en liten del av kostnaderna för privat tandvård.
Vissa kommuner ordnar förberedande undervisning före den grundläggande utbildningen för elever som ännu inte har tillräckligt bra språkkunskaper för den vanliga undervisningen.
På servicestället hjälper FPA:s och Skatteförvaltningens experter invandrare som kommer till Finland för att arbeta i frågor som rör beskattning och social trygghet.
Tfn: (09) 8392 4682
Tjänsten ger dig förslag på olika kollektivtrafikförbindelser från ett ställe till ett annat.
Anställningsrådgivningen har öppet på tisdagar och onsdagar klockan 9–11 och 12–15.
I Finland erbjuder kommunerna tjänster för bostadslösa.
Beskriv dina arbetsuppgifter och de färdigheter som du lärt dig i arbetet.
Du kan omfattas av den finländska sociala tryggheten endera på basis av stadigvarande bosättning eller på basis av arbete.
Läs mer: Bibliotek.
Resplan för cycling och gångfinska _ svenska _ engelska _ ryska
Vid kommunalval och Europaparlamentsval har dock också andra länders medborgare som bor i Finland rösträtt.
Du bör observera att den partiella förtida ålderspensionen permanent minskar beloppet på den slutliga ålderspensionen.
Dessutom finns det gym av flera olika slag.
Ditt betyg, inträdesprovet och din arbetserfarenhet kan påverka antagningen.
Du ska besöka beskickningen eller tjänstestället inom tre månader efter att ha gjort ansökan på internet.
I Finland utkommer även den ryskspråkiga tidskriften Spektr.
Fråga mer på din mottagningscentral.
Kommunerna ordnar förskoleundervisning.
Grundskolan består av lågstadiet (alakoulu) och högstadiet (yläkoulu).
Graviditetspreventionfinska
Information om kyrkans familjerådgivningfinska _ svenska
Det är bra att diskutera bytet av efternamn även med barn som ännu inte har fyllt tolv år.
Om du flyttar permanent från Finland eller vistas utomlands två år utan avbrott återkallas ditt uppehållstillstånd.
Utred din situation tillsammans med socialarbetaren: hur mycket kan du betala i hyra, och kan du få hyresstöd.
Stöd för alkoholisterfinska _ svenska _ engelska
Privata hälsovårdstjänster
linkkiEsbo stad:
Hälsovård för anställda och företagare
När du flyttar till Finland måste du göra en flyttanmälan och gå och registrera dig vid magistraten (maistraatti) på din egen hemort.
Försäkringen får inte vara en vanlig reseförsäkring.
Arbets- och näringsministeriet svarar för beredningen av ärenden i anslutning till integrationen av invandrare i Finland.
du har en fast anställning eller motsvarande avtal för ett arbete som du utför i Finland
Du kan ansöka om invaliditetspension med en blankett som du får från FPA.Som bilaga till ansökan krävs B-utlåtande av läkare.
Social kreditgivning
Läs mer om finska medborgares rättigheter och skyldigheter på InfoFinlands sida Finskt medborgarskap.
Civilvigsel kan enligt lag förrättas av en häradsskrivare som arbetar vid magistraten (maistraatti) eller en lagman eller tingsdomare som arbetar i tingsrätten (käräjäoikeus).
Detta är särskilt viktigt om du upptäcker att det samlas vattenånga eller fukt på fönstren när du lagar mat.
stadfäster lagarna,
Vem är flykting?
När du fyllt i ansökningen i tjänsten har du tre månader på dig att styrka din identitet.
Mariegatan 28, 67200 Karleby
Till exempel studerande vid den samhällsvetenskapliga eller den humanistiska fakulteten utexamineras inte nödvändigtvis till ett yrke.
Du kan lära dig att spela ett instrument, sjunga i kör, gå på konserter och festivaler eller till och med sjunga karaoke.
Patientombudsmannens verksamhetfinska _ svenska _ engelska
Läs mer: Registrering som invånare, Hemkommun i Finland.
Domstolen undersöker inte varför man ansöker om skilsmässa.
Förlossningarfinska _ svenska
Finnvera är ett specialfinansieringsbolag som ägs av finska staten.
Stöd för närståendevårdfinska _ svenska
Gymnasium
Ungdomar under 15 år bestraffas inte för brott.
linkkiRovaniemi stads ungdomstjänster: Hyresbostäder i Rovaniemifinska
Dessutom erbjuds åldringar i Esbo egna tjänster, till exempel hemvårdens tjänster.
Tfn 09 819 55360
Om barnet dessutom behöver avgiftsbelagd småbarnspedagogisk verksamhet arrangeras denna på samma ställe som förskoleundervisningen, dock med undantag för skiftesvård.
Socialarbetare 016-322 3088, 040-576 8914
Om du har finska nätbankskoder kan du även köpa personligt resekort på HRT:s webbplats.
En sådan stödperson kallas doula.
Även i museikvarterens övriga byggnader finns utställningar om stadens kulturhistoria och utställningar med ITE-konst.
NEJ: PVC-förpackningar med märkningen 03, förpackningar som innehåller rester av farliga ämnen såsom målarfärg eller kemikalier, plastföremål, leksaker, tandborstar, vattenkannor och så vidare
Om du inte betalar räkningen eller kommer överens om en betalningsplan kan skulden slutligen gå till utmätning (ulosotto).
Det ger lån till nya företag och redan aktiva företag.
Vid behov förs barnet till stadens hälsostation.
Efter det första året kallas man till barnrådgivningen ännu minst sex gånger.
Familjerådgivningar finns på många orter.
Om barnet får medborgarskap i ett EU-land, ska du ansöka om registrering av EU-medborgares uppehållsrätt för barnet i Migrationsverkets e-tjänst Enter Finland eller vid Migrationsverkets serviceställe.
Handikapporganisationer i Finlandfinska _ svenska
upprättande av stadgar
En utredning över att du har tillräckliga medel för din försörjning i Finland.
Om bara en av parterna står som köpare är denne ägare till egendomen när samboförhållandet upphör.
Du kan ansöka om stipendier hos olika stiftelser (säätiö).
Nationellt hjälpsystem till offer för människohandel i Finland
Du måste dock själv skaffa gymnasieböckerna.
I tjänsten Reseplaneraren (Reittiopas-palvelu) kan du söka information om kollektivtrafikens rutter i huvudstadsregionen.
En person som står under förmynderskap klarar inte av att sköta sina angelägenheter utan de sköts av en intressebevakare.
TE-byrån eller kommunen anvisar dig vid behov till integrationsutbildning.
Hemförsäkringen ersätter till exempel skador på möbler och andra ägodelar.
Tidsbeställning till tillståndstjänstenfinska _ svenska _ engelska _ samiska
Flexibel och partiell vårdpenning
Du hittar mer information om den offentliga hälso- och sjukvården på InfoFinlands sida Hälsovårdstjänster i Finland.
Hälsostationernafinska _ svenska
ett löneintyg för de senaste sex månaderna om dina inkomster har ökat.
Inom två veckor efter att barnets födelse registrerats skickar magistraten en blankett hem till modern.
En asylsökande är alltså inte en flykting (pakolainen).
Polisen kan utfärda identitetskort för en utlänning som
Läs mer på InfoFinlands sida Samboförhållande.
Meddela namnet till magistraten.
Om du inte är stadigvarande bosatt i Finland
Pålitlighet och att hålla tidtabeller
Många skolor håller kontakt med föräldrarna med hjälp av webbtjänster.
du inte söker ett jobb som TE-byrån föreslår för dig
du inte tar emot ett jobb som erbjuds till dig
På många orter finns medborgarinstitut, som kommunerna upprätthåller.
Hörselskadade
Den sociala tryggheten i Finland
Ansökan om uppehållstillstånd är avgiftsbelagd.
Du kan även besöka servicestället In To Finland i Kampen i Helsingfors för att fråga om beskattningen.
Vad ska jag beakta när jag använder bastun i min bostad?
Besöksadress: Ämbetshuset, Torggatan 40, 67100 Karleby
Mer information om graviditet och förlossning hittar du på Vanda stads mödra- och barnrådgivning på Internet (Nettineuvola).
Läs mer på InfoFinlands sida Utländska examina i Finland.
Du hittar kontaktuppgifterna vid din församling.
Arbetsgivare behöver inte ge dig ett arbetsintyg på eget bevåg.
grundtryggheten för arbetslösa
Upphovsmannen som deltar i tävlingen överlåter rätten att kopiera verket och ändra verkets format och storlek i den omfattning som krävs för att visa verket.
Ett tidsbestämt avtal (Määräaikainen vuokrasopimus) innebär att hyresvärden och hyresgästen från början kommer överens om när avtalet upphör.
Lönejämförelse finska _ engelska
När du väntar barn
Information om brottfinska _ svenska _ engelska
Det finns bostadsrättsbostäder i de största kommunerna.
Bibliotekfinska _ svenska _ engelska
Stöd och verksamhet för flickorfinska
Stipendiet kan täcka hela läsårsavgiften eller en del av den.
Också borgerliga vigslar förrättas på magistraten.
Läs mer på InfoFinlands sida Abort.
du återkallar din asylansökan
I Finland förväntar människorna sig att man verkligen menar det man säger.
I Finlands talas tre olika varieteter av samiska.
Invandrarenheten hjälper också personer som fallit offer för människohandel.
Då klär barn sig ut till häxor och går runt i grannskapet för att dela ut videkvistar som de dekorerat.
Idrottsklubbarfinska
Skolhälsovårdfinska _ svenska _ engelska
Eldstadstorget 1 eller Kopparbergsvägen 10 B, vån.
Förlovningen är frivillig och krävs inte i lag.
Du kan gå till en privat läkarstation även om du inte har rätt att använda den offentliga hälso- och sjukvården i Finland.
I Karleby finns en ortodox kyrka.
I Finland kan makarna byta efternamn när de gifter sig.
Lämna inte linor eller annat fiskeavfall i naturen.
Frivillig återflyttningfinska _ svenska _ engelska
Vid MoniNet kan du få information om hobbyer, till exempel kurserna vid medborgarinstituten eller föreningsverksamhet.
Hurdant utkomstskydd för arbetslösa får företagare i Finland?
mån–fre kl. 8.00–16.00 (för personligt möte måste du boka tid)
de partier som har minst en riksdagsledamot,
Tjänsten Internationell personbeskattning tillhandahåller information om beskattningen av inkomster från utlandet och beskattningen av arbete utomlands samt hur en flytt utomlands påverkar beskattningen.
Unga kan prata om sina problem med hälsovårdaren på den egna skolan eller läroanstalten.
För att få vård måste du ha ett europeiskt sjukvårdskort.
Om du vill söka en av stadens hyresbostäder ska du fylla i en ansökningsblankett för hyresbostäder.
Efter studierna på andra stadiet kan du gå vidare till högskoleutbildning.
linkkiTrafiksäkerhetsverket:
Ingången till byrån för ungdomstjänster ligger på torgsidan. Ta trappan upp till andra våningen.
Bioavfall komposteras till mylla.
Läs mer: Barns hälsa.
I vissa kommuner har barnet rätt till småbarnspedagogik på heltid även då den ena föräldern är hemma.
I Helsingfors finns även privata daghem vars verksamhetsspråk är engelska, ryska, tyska, franska eller spanska.
Rådgivning ges både per telefon och via e-post:
Om du omfattas av den finländska sociala tryggheten kan du ansöka om arbetslöshetsstöd.
Evenemangfinska _ svenska _ engelska _ ryska _ kinesiska
Gemensam ansökan till yrkeshögskolorfinska _ svenska
När du tar med dig en bil till Finland som flyttsak, måste du tullanmäla den.
Betjäning ges på finska och svenska samt i mån av möjlighet även på engelska.
Servicepunkt för socialarbete och socialhandledningfinska
Läs mer på InfoFinlands sida Arbetarskydd.
Kontaktuppgifterna till rådgivningsbyråerna hittar du på Vanda webbplats.
Du kan fråga om doulaverksamheten på din hemort vid rådgivningen.
Många skaffar sig en julgran som pyntas.
Till Kalkkers kan du även komma utan uppehållstillstånd.
Visumbehovet till Schengenområdet och av
Upprätthåll ditt kunnande, följ aktuella händelser och nyheter i din bransch, delta i kompletteringsutbildning och utveckla tidigare kunskaper.
Om du har frågor kring stödtjänsterna för äldre, kontakta Esbo stads rådgivning för seniorer.
De flesta invånarna är finskspråkiga.
Storgatan 3, 67100 Karleby
Då är den inte nödvändigtvis mycket dyrare än den kommunala småbarnspedagogiken.
Läs mer: Problem med uppehållstillstånd.
Kela betalar stödet direkt till skötaren eller dagvårdsproducenten.
Vid Helsingfors vuxengymnasium finns en linje avsedd för invandrare över 17 år, där du kan avlägga hela eller en del av den grundläggande utbildningen.
Man kan också söka skilsmässa ensam.
Du måste skriva alla prov på högst tre efter varandra följande examenstillfällen.
Bokning av tid till barnatillsynsmannen:
Du kan också ansöka om personbeteckning från magistraten.
Ledd motion kan vara till exempel jympa eller promenader, löpning eller skidåkning i grupp.
I förskoleundervisningen skaffar sig barnet förberedande färdigheter inför grundskolan.
du studerar i Finland och dina studier räcker minst två år
Du behöver ha minst 560 euro disponibla medel i månaden för att kunna betala för boende, mat och andra utgifter.
Om du är intresserad av att grunda ett eget företag, gå in på InfoFinlands sida Att grunda ett företag.
Tfn (09) 4711
Mer information om brottsanmälan hittar du på InfoFinlands sida Brott.
EU-medborgare som är i det finska rösträttsregistret kan också ställa upp som kandidat i Finlands Europaparlamentsval.
På Furumo begravningsplats finns även ett gravområde för konfessionslösa. Där kan de avlidna begravas som inte hörde till ett religionssamfund.
Religionsundervisning måste ordnas när det finns minst tre barn som bekänner en viss religion i kommunen.
Tolken ska vara myndig, så egna minderåriga barn kan inte användas som tolk.
Kom ihåg att returnera eller förnya dina lån i tid.
Arbetstagarförbunden är organiserade under tre centralförbund för löntagare.
Kalkkers håller öppet kl. 22–6.
Om magistraten registrerar din uppehållsrätt, registreras dina personuppgifter automatiskt även i befolkningsdatasystemet.
en utländsk examen, som ger möjlighet till universitetsstudier i det land där du avlagt examen
har fyllt 18 år och
Ungdomscentralen Nuppi (nuortenkeskus Nuppi) hjälper ungdomar med missbruksproblem, Internetberoende eller spelberoende.
För alltid farligt avfall till insamlingsställe.
p. 050-593 0165
Om du behöver omedelbar krishjälp, kan du också ta kontakt med social- och krisjouren.
Ett efternamn som maken eller makan har fått från sitt tidigare äktenskap kan inte väljas som efternamn.
I Rovaniemi finns mångsidiga motionsmöjligheter.
Tfn (09) 839 21064
Flick- eller pojkvän till en finsk medborgarefinska _ svenska _ engelska
Våren 1918 befann sig Finland i inbördeskrig som kämpades mellan de röda gardena som representerade arbetarna och de vita skyddskårerna som representerade borgarna och markägarna.
Mer information om tjänster för handikappade får du från Mellersta Österbottens social- och hälsovårdssamkommun Soites handikapptjänster per telefon: 040 804 2122.
Lapplands centralsjukhus
På InfoFinlands sida EU-medborgare hittar du information om flytt till Finland av andra skäl än som asylsökande.
Kort vistelse i Finland
I Finland är vissa yrken reglerade.
Barn under 17 år kallas till tandkliniken för undersökning med cirka två års mellanrum.
Eftersom Finland lyckades försvara sitt territorium i krigen kort efter att landet hade blivit självständigt har krigen under 1900-talet betraktats som den tid då Finlands självständighet etablerades.
Du kan även ändra kontaktspråket senare.
Om du misstänker att du blivit utsatt för diskriminering då du sökt arbete eller på arbetsplatsen ska du först ta upp detta på din arbetsplats.
linkkiFörbundet för ungdomsbostäder rf:
Registrering av uppehållsrätten för EU-medborgare sker inte per automatik.
Information om krissituationer och sorgfinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Upphovsrätt:
Yrkesutbildningfinska _ engelska
Man försöker alltid ingripa i problem redan innan de blivit alltför stora.
Handläggning av ansökan om uppehållskort är avgiftsbelagd.
lägre eller högre högskoleexamen vid universitet eller högskola
Studierna är allmänbildande.
I skolan arbetar även en psykolog eller en kurator.
tillhörighet till en viss grupp i samhället eller
God natt!
den regelbundna arbetstiden
I Finland anses det vara välartat att ta hänsyn till och lyssna på andra.
A1 – ASE 1
Val av gren och grupp
Ett tillstånd av hyresvärden behövs alltid för detta.
Arbetsgivaren ska välja den sökande som har de bästa meriterna för uppgiften.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
anstaltsvård
Om en företagare blir sjuk
Hjälptelefonfinska _ svenska _ engelska
Ett tidsbestämt hyresavtal upphör automatiskt utan uppsägning på den dag som antecknats i avtalet.
Åldershörselfinska
På InfoFinlands sida Vad är en familj?
I Finland bor många människor i hyresbostäder.
Ett bevis på stadigt sällskapande kan till exempel vara att er avsikt är att ingå äktenskap i Finland.
Förberedande för yrkesutbildning
Om du inte är kund hos arbets- och näringsbyrån görs den inledande kartläggningen och integrationsplanen på socialbyrån.
Du kan få arbetslöshetsersättning tidigast från den dag då du gjort anmälan vid TE-byrån.
Mer information om personbeteckningen hittar du på InfoFinlands sida Registrering som invånare.
Sjukdagpenning betalas för högst 300 vardagar.
rehabiliteringskurser för personer med en viss sjukdom
pengar
till ett gott bemötande: patientens människovärde, övertygelse och integritet ska respekteras
Syftet med tjänsterna är att hjälpa den handikappade att vara delaktig i samhället och underlätta livet med handikappet.
Kontaktuppgifter till magistratfinska _ svenska _ engelska
och integrationsplanen tillsammans med dig om du anmäler dig till TE-byrån som arbetslös arbetssökande.
Försörjningsförutsättning för make/maka till en finsk medborgare
De finns runtom i huvudstadsregionen.
Information om erkännande av examen för yrken inom hälsovårdenfinska _ svenska _ engelska
Du har inte lämnat till exempel skatter, böter, underhållsbidrag eller sjukhusavgifter obetalda.
Under vårdledigheten kan du ansöka om hemvårdsstöd av Fpa.
Du kan ansluta dig till fackförbundet i din egen bransch.
Social- och krisjouren 24 h
linkkietsilaakari.fi:
Lätt motion kan även vara till exempel trädgårdsskötsel, städning eller snöskottande, d.v.s. så kallad vardagsmotion (hyötyliikunta).
linkkiKarleby evangelisk-lutherska församlingssammansutning:
Senioruniversitetet ordnar föreläsningsserier, kurser och studieresor.
I Finland är det vanligt att kvinnor arbetar, även om de har barn.
Handikappbidrag för vuxna betalas till 16–64-åringar.
Du kan också söka information om privata jurister på till exempel Finlands Juristförbunds (Suomen Asianajajaliitto) webbplats.
Helsingfors har cirka 650 000 invånare. 78 procent av invånarna har finska och 6 procent har svenska som modersmål.
Om du inte har ett jobb eller om du blir arbetslös, anmäl dig på arbets- och näringsbyrån senast på din första dag som arbetslös.
Denna person ansvarar i sista hand för att de tillstånd som krävs för att göra videoklippet skaffas, att tillstånden är vederbörliga, att eventuellt material i videoklippet som en tredje part har upphovsrätt till används vederbörligt samt för eventuella upphovsrättsavgifter och upphovsrättsliga krav.
I Finland kan man avlägga högskolestudier både vid yrkeshögskolor och vid universitet.
Vissa stipendier kan även täcka andra kostnader.
Underhållsstöd
FPA kontaktuppgifterfinska _ svenska _ engelska
Strykjärnet ska också kopplas loss från vägguttaget.
en kopia av överenskommelsen mellan dig och din arbetsgivare om att du under en viss tid ska arbeta på deltid.
Fråga mer vid rådgivningstjänsterna för invandrare, utbildningsväsendet i din hemkommun eller studievägledarna vid lokala läroanstalter.
Vanligtvis när du söker ett jobb, skickar du en jobbansökan och ditt CV, alltså din meritförteckning, till arbetsgivaren.
Ledd motion ordnas till exempel av kommuner och idrottsklubbar.
Vissa länder har också konsulat i andra städer.
Låt alltid barnets intressen gå först när ni fattar beslut.
Om makarna har upprättat ett äktenskapsförord delas egendomen vid skilsmässa eller när den ena makan avlider i enlighet med det. Om makarna har upprättat ett äktenskapsförord delas egendomen i enlighet med det.
Branschförbunden är intressebevakningsorganisationer för företag i olika branscher.
Då var södra Esbo fortfarande hav.
Om du är sjuk under en längre tid får du vanligtvis först under ungefär ett års tid sjukdagpenning.
Du kan även publicera en egen annons.
Uppehållstillstånd för företagarefinska _ svenska _ engelska
Lånet återbetalas det vill säga amorteras en gång i månaden.
Läs mer på Vanda stads webbplats.
Det bör finnas en brandvarnare på varje våning.
När du behöver rehabilitering behöver du först ett läkarutlåtande.
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
Dessa tjänster är avsedda för människor som har en hemkommun i Finland.
Du kan också ansöka om ditt första visum i Finland, om din familjemedlem är finsk medborgare och du själv är medborgare i ett visumfritt land, det vill säga du inte behöver visum för att komma till Finland.
Planerar du att flytta från Finland till ett annat land?
Om du har ett bostadslån i en utländsk bank, ska du själv ge uppgifterna om lånet till skattemyndigheten.
Läs mer på InfoFinlands sida Stöd till gravida och Stöd efter barnets födelse.
Läs mer:
Penningunderstöd för utländska forskarefinska _ engelska
Social trygghet för dig som flyttar till Finland(pdf, 560 kb)finska _ svenska _ engelska _ ryska _ estniska
Jämför elpriserfinska
linkkiEsbo församlingar:
Mental hälsafinska _ svenska
Enligt Finlands lag är alla barn jämställda oavsett bakgrund eller ålder.
Om den unga inte är trygg i sitt eget hem, kan hen kontakta Finlands Röda Kors De ungas skyddshus.
Sökning av ägarbostäderfinska
Privatpersoner lägger även ut tidningsannonser om bostäder som de hyr ut.
linkki4V:
Jag misstänker att jag har blivit diskriminerad när jag letade efter bostad.
Väestöliittos mångkulturella arbete stödjer invandrafamiljer.
Också äldre människor har nytta av att röra på sig, eftersom motion upprätthåller den fysiska konditionen och funktionsförmågan.
studerande
Det gäller även arbetstagare som blivit utsända utomlands av sin finska arbetsgivare.
Kamrersvägen 2 A, vån. 4
Också förlossningen blir lättare.
Friluftsliv och vandring
När en gift kvinna får ett barn registreras kvinnans make automatiskt som barnets far i befolkningsregistret.
Information om studier i Finland hittar du på InfoFinlands sida Utbildning.
Du kan få uppehållstillstånd på grund av familjeband om ditt barn bor i Finland.
Arbetsgivaren ska teckna en olycksfallsförsäkring (tapaturmavakuutus) åt sina anställda.
tfn 016 322 2269
En integrationsplan utarbetas för dig åtminstone om
Privata dagvårdsplatser söks direkt på daghemmet.
Problem i äktenskap eller parförhållande
I Karleby ges gymnasieutbildning för ungdomar vid Karleby finska gymnasium och Karleby svenska gymnasium, samt för vuxna vid Karleby vuxengymnasium.
Varje anställd har rätt till ett jämlikt och icke-diskriminerande bemötande när de söker jobb och på arbetsplatsen.
På vintern är många motionsslingor skidspår.
Du väljer själv hur mycket studielån du vill ta.
Gymnasiet kan också avläggas på två eller fyra år.
Lyssna på finska dialekterfinska
Du kan ringa skyddshuset under alla tider på dygnet.
Fristående examen (näyttötutkinto) är ett sätt att bevisa sin yrkeskunnighet.
Stadens hyresbostäder är ofta billigare än bostäder som man hyr av företag eller privatpersoner.
skött bostaden omsorgsfullt och
Esbo social- och krisjour vid Jorv sjukhus betjänar personer som bor i Grankulla.
Information om att arbeta och driva ett företag i den europeiska unionenfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
Om du är intresserad av att grunda ett eget företag, gå in på InfoFinlands sida Att grunda ett företag.
Om du behöver psykiatrisk vård kan du kontakta din hälsocentral.
linkkiFinnkino:
Om du omfattas av den sociala tryggheten i Finland kan du ansöka om bostadsbidrag för boendekostnader hos FPA.
Hemförsäkringar säljs av många försäkringsbolag i Finland.
Om du är minderårig och vill göra abort behöver du inte tillstånd av dina föräldrar.
Parker för invånare och öppna daghemfinska _ svenska _ engelska
Ansök om tillståndet i ditt hemland eller i ett annat land där du vistas lagligt. Du kan också ansöka om ditt första uppehållstillstånd i Finland om din make eller maka är finsk medborgare och du själv är medborgare i ett visumfritt land, det vill säga du inte behöver visum för att komma till Finland.
Arbetsgivaren är också skyldig att sörja för arbetstagarnas säkerhet och hälsa i arbetet.
Avfallshantering och återvinning
Du kan skriva till Väestöliitto på dari, kurdiska (sorani), persiska, finska, ryska, engelska eller svenska.
Behöver du juristhjälp? Barns och ungas problem
Inledande kartläggningfinska _ engelska
De öppna universiteten tillhandahåller universitetskurser.
behovsprövad rehabilitering
Kassen eller påsen får vara högst 30 l stor.
Företagarens företagshälsovård (työterveyshuolto)
Motionsmöjligheterfinska
Om du behöver råd i sådant som rör fostran av barn eller barns utveckling, kan du boka en tid hos familjerådgivningen (perheneuvola).
Att grunda ett företag
Du får information om hälsovårdstjänster i Finland på InfoFinlands sida Hälsa.
Om din lön uppgår till minst 696,60 € i månaden, har du rätt till de flesta av FPA:s förmåner.
Skyddshuset har öppet kl. 17–10, telefonjouren betjänar dygnet runt.
Det är dessutom möjligt att studera vid den öppna yrkeshögskolan.
Fråga närmare av FPA.
eBiblioteketfinska _ svenska _ engelska
Pensionsskyddscentralen sköter centraliserat frågor som rör pensionsskyddet.
Ta med dig ett identitetsbevis och ansökningsbilagorna i original.
Det innebär att du inte behöver betala för de hjälpmedel som du behöver för att klara dig i vardagen.
Om du använder andra fiskeredskap ska du ha ett fisketillstånd.
tullen,
Begravningsbidrag
Statens lokalförvaltning
Tfn 09 7562 2260
När du har bokat en telefontid, ringer FPA:s servicerådgivare upp dig vid överenskommen tidpunkt.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
I Finland omfattas högskolestuderande av studerandehälsovården.
Tolken har sekretessplikt och får inte berätta inte om dina angelägenheter för andra.
Cykling
Föräldrarnas uppehållstillstånd kan dock påverka vilka stöd familjen kan få.
från vilket land du flyttar till Finland.
Du kan köpa kondomer i affärer, på bensinstationer, kiosker och apotek.
Det är bra att gå på läkarundersökning första gången före utgången av den fjärde graviditetsmånaden.
Du kan sättas i karens till exempel om:
till att patientens modersmål och kultur beaktas i den mån det är möjligt
Ansök om dagvårdsplats på Internet.
Bouppteckning
Både kvinnan och mannen har rätt att söka skilsmässa.
En del av kurserna är avsedda för personer som ska starta eget företag och en del för dem som redan har eget företag.
Arbetsplatser vid stadenfinska _ svenska _ engelska
Tfn (09) 816 30300
Tjänster för handikappade är till exempel personlig assistans, serviceboende, färdtjänst och ombyggnadsarbeten i bostaden.
Nödcentraloperatören ser var du är, när du ringer ett nödsamtal via appen.
En sjukskötare eller läkare besvarar ditt samtal.
På dessa sidor redogörs det för hurdant ekonomiskt stöd barnfamiljer kan få i Finland.
De ordnar föräldramöten och berättar för föräldrarna om barnets studier.
Sexuellt våld är alltid ett brott, även i äktenskap.
linkkiTidningarnas föbund:
Förvaltningsdomstolen kan antingen avslå besvären eller sända ärendet till Migrationsverket för ny behandling.
Alla barn som har sitt stadigvarande boende i Finland har läroplikt, vilket innebär att de måste delta i den grundläggande utbildningen.
På InfoFinlands sida Flykting hittar du mer information avsedd för flyktingar.
Läs mer på InfoFinlands sida Pension.
Barnet lär sig också olika färdigheter som hjälper hen att lära sig ytterligare nya saker.
_ tjeckiska
Om du använder en egen bil ska du enligt lagen ha en trafikförsäkring.
linkkiEsbo vuxengymnasium Omnia:
De olika språkversionerna av InfoFinlands är identiska.
El
Om du har fått ditt första barn kan stödpersonen ofta även tillbringa nätterna på sjukhuset.
Miehen Linja är en tjänst för invandrarmän som har utövat våld eller fruktar att de kommer att utöva våld mot sin maka eller någon annan familjemedlem.
Båda språken har långa traditioner i Finland.
Undervisningsutbudet varierar från år till år, så det lönar sig att kontrollera aktuella kurser på institutets webbplats.
Under denna tid kan du inte resa utomlands.
Stora midsommareldar hör till de finländska midsommartraditionerna.
Genom läroavtalsutbildning (oppisopimuskoulutus) (ungdomar och vuxenstuderande)
Gör hyresavtalet alltid skriftligt.
Information om Helsingforsfinska _ svenska _ engelska
Den finansieras med skattemedel och är därför kostnadsfri för familjerna.
Stöd för vård av barn i hemmet.
1948 VSB-avtalet mellan Finland och Sovjetunionen
sambor
Uppehållstillstånd
Du kan söka teaterföreställningar i evenemangskalendrarna på sidorna myhelsinki.fi och stadissa.fi.
Ungdomsgårdenfinska _ svenska _ engelska
Varje religiöst samfund bestämmer själv vilka villkor som gäller för vigseln och hurudan vigselceremonin är.
Du kan även ansöka om uppehållstillstånd på någon annan grund.
Om det behövs kan du också anlita en tolk.
De flesta arbetsgivare värdesätter att den anställda vill utveckla sig i sitt arbete och inhämta nya kunskaper.
Vuxna kan avlägga gymnasiestudier på vuxengymnasiet.
Kontrollera också om du till exempel har rätt till bostadsbidrag eller utkomststöd.
För att du ska kunna få ett bostadslån måste du ha tillräckliga inkomster för att betala tillbaka lånet utan problem.
följa de överenskomna arbetstiderna
Du behöver inte alltid boka tid för att besöka TE-byrån.
Läs mer på sidan: Skattedeklaration och beskattningsbeslut.
Du kan inte få hemvårdsstöd om barnet går i den kommunala dagvården.
Ordföljden är friare än i många andra språk.
Läs mer på InfoFinlands sida Familjeledighet.
Akademiskt erkännande av examina betyder
Nybörjarkurs i finska, Tavataan taasengelska _ franska _ tyska _ bulgariska
Vårdnadsavtalet ingås antingen på rådgivningsbyrån före barnets födelse eller hos barnatillsyningsmannen efter barnets födelse.
När du ställt ansökan ska du besöka Finlands beskickning närmast dig för att styrka din identitet och visa upp originalexemplaren av ansökningsbilagorna.
Inledande kartläggning
I Finland betalas skatt på pensionerna.
Daghem som ger förskoleundervisningfinska _ svenska _ engelska
Krisen kan till exempel ha med våld, parförhållandet eller barnens problem att göra.
Vid posttraumatiskt stressyndrom väcker olika situationer minnesbilderna från den traumatiska situationen, vilket orsakar kraftig ångest.
Kravet på tillräcklig inkomst tillämpas dock inte på föräldern om barnet fötts innan föräldern anlänt till Finland och föräldern har flyktingstatus i Finland.
På Omnia kan man studera många olika yrken.
Du kan ansöka om tillståndet på internet via tjänsten Enter Finland.
Om du har problem eller oklarheter med uppehållstillståndet, kan du ta kontakt med migrationsverket.
Annan allmän information i ämnet finns på InfoFinland-sidan Flytta till Finland.
Man kan också bo korta tider i en anstalt.
Om du har omskurits (ympärileikkaus) innan du kom till Finland öppnas din slidmynning med operation (avausleikkaus) i samband med förlossningen.
Du får samtidigt även en finsk personbeteckning.
egendom
Mottagare av statsförvaltningens språkexamina, svenska språketfinska _ svenska
du inte har en ägarbostad på samma område; och
Helsingfors evenemangskalenderfinska _ svenska _ engelska
Du kan också vara partiellt vårdledig.
linkkiFinlands Advokatförbund:
Sidunderhåll
I Finland är försvarandet av familjens eller släktens heder inte en godtagbar anledning till hot, påtryckningar eller våld.
Grundläggande utbildning
Information om stiftelser och penningunderstödfinska _ svenska _ engelska
linkkiHelsingforsnejdens kontakttolkcentral:
Barnets föräldrar eller vårdnadshavare kan inte vägra vård om barnet behöver den.
Läs mer: Brott.
Kontrollera vad hyresavtalet säger till exempel om villkoren för hyresförhållandet och om uppsägningstiden.
Du kan läsa mer om värderingar och seder i det finländska samhället på sidan Finländska seder.
Till exempel i Lappland äts mycket renkött, medan man i kustregionerna äter fisk.
Du kan också sluta arbeta.
Ta med dig ett giltigt ID-kort eller pass.
Resekortet gäller i lokaltrafikens bussar, närtågen, metron, spårvagnarna och Sveaborgsfärjorna.
Arbetshälsa och rekreation
På biblioteket kan det även finnas sagotimmar och spel för barn.
Vi ger stöd och råd åt invandrarkvinnor som blivit utsatt för våld eller lever under hot om våld.
Där är det ingen som frågar om du har uppehållstillstånd.
Om du måste sköta ärenden med finländska myndigheter, men inte kan finska eller svenska och det inte heller finns något annat språk som både du och myndigheten talar, kan du i vissa fall ha rätt till tolkning.
Rovaniemi stads familjerådgivning
Varken du eller din partner får vara gift med någon annan.
Evenemangfinska _ svenska _ engelska _ ryska
I tjänsten medverkar Helsingfors-info, magistraten i Nyland, skatteförvaltningens och FPA:s tjänst In To Finland, NTM-centralen i Nyland, Pensionsskyddscentralen och Helsingforsregionens handelskammare.
Mer information om hurdana kunskaper de olika nivåerna avser i praktiken får du på Utbildningsstyrelsens (Opetushallitus) webbplats.
en kopia av hyresavtalet och en utredning över hyresbeloppet (hyresbostad)
Om du är medborgare i ett annat land måste du besöka arbets- och näringsbyrån.
tfn. 09 6850 120
På InfoFinlands sida Fostran av barn i Finland finns information om hur barn fostras i Finland.
Läs mer: Bibliotek.
Om du får avslag på din ansökan om uppehållstillstånd eller om förvaltningsrätten avslår ditt överklagande, måste du lämna Finland.
Midsommar är en högtid som firas nära sommarsolståndet.
Tjänsterna är avgiftsfria.
Innan du kan ansöka om uppehållstillstånd måste du skaffa dig en studieplats i Finland.
Arbets- och näringsbyråeran upprättar även integrationsplaner för invandrare som är klienter vid arbets- och näringsbyrån.
Om hen försöker göra detta kan du polisanmäla hen.
Bostadsbidrag beviljas för skäliga boendekostnader.
Vanligtvis är barnets mor eller far vårdnadshavare.
Du kan även göra det personligen på Migrationsverkets tjänsteställe.
Nollalinja är avsedd för både kvinnor och män.
Muslimerna i Helsingfors har sitt eget gravkvarter på Furumo begravningsplats i Vanda.
Barnet kan få uppehållstillstånd på grund av familjeband om hans/hennes föräldrar har uppehållstillstånd i Finland och en förälder bor i Finland.
Till exempel föräldrarna får inte tvinga sitt barn att gifta sig.
Du kan ta upp problemet med proffs inom hälsovården eller företagshälsovården, som kan slussa dig vidare i vårdsystemet, eller direkt kontakta Soites missbrukstjänster, tfn 040 8068 101.
Jämställdhet i arbetslivet
Som asylsökande har du rätt att använda ett rättsbiträde under samtalet.
Vissa betalningar går emellertid direkt till utmätning.
FPA beställer tolken.
Utbildning på andra stadiet
Kontaktuppgifter till kontorenfinska _ svenska _ engelska
Ansökan om progressiv inkomstbeskattningfinska _ svenska _ engelska
Karleby har satsat på att förbättra förhållandena för cyklister.
Det är artigt att ta av sig skorna när du går in i någons hem.
MoniNet
Broschyr om erkännande av examen(pdf, 102,14 kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ kinesiska _ persiska _ arabiska
Lönen och utbetalning av lönen
Valtakatu 16
Läs mer: Universitet och Yrkeshögskolor.
Du kan ansöka om stödet vid socialbyrån i din egen kommun.
linkkiEdupoli:
Högskoleutbildningfinska
Hjälp vid ekonomiska problem
Grundläggande utbildning.
Du får blanketten hos arbetskraftsmyndigheten i ditt hemland.
I nödfall får du vård inom den offentliga hälso- och sjukvården fastän du inte har en hemkommun i Finland eller rätt till vård på grund av arbete.
Vinnaren belönas med en tabletdator.
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
Jag upplever att jag blir osakligt bemött på min arbetsplats.
Arbetsgivaren får inte diskriminera de anställda när han eller hon fattar beslut om fördelning av arbetsuppgifter, erbjudande av möjligheter till avancemang eller upphävande av anställningen.
På det finska utrikesministeriets webbplats finns en förteckning över andra länders beskickningar i Finland.
Anmälan till grundskolan sker vid den skola som anges i ett brev som varje ny elev får hem eller per telefon till skolan.
som har ifrågavarande kommun som hemkommun och
Tfn (09) 310 6611 / 116 117
Under tiden kärnkraftverket uppförs kommer som mest upp till 3 000–4 000 personer att arbeta på området.
Telefonnumret är 09 471 71110.
Om kristna fester kan du läsa mer på webbplatsen för evangelisk-lutherska kyrkan i Finland.
Familjemedlem till en person bosatt i Finland
På vissa arbetsplatser måste man kunna både finska och svenska.
Underhållsbidragets belopp beräknas utifrån barnets underhållsbehov och föräldrarnas underhållsförmåga.
Musikfestivaler är populära, särskilt på sommaren.
Föräldradagpenningar är skattepliktiga inkomster och följaktligen behöver du ett skattekort (verokortti).
Om du inte har en hemkommun i Finland eller om du inte omfattas av sjukförsäkringen i Finland, kan du ändå ha rätt till vård eller ersättningar från FPA på någon annan grund.
praktik
Att enbart använda bostaden för det avsedda ändamålet.
Make/maka till en utländsk medborgare
Offentliga hälso- och sjukvårdstjänster samt socialtjänster är kommunernas ansvar i Finland.
18–22 år och har bott i Finland i flera år
Du kan ringa nödnumret gratis från alla telefoner.
Man kan också vända sig till förtroendemannen till exempel med frågor om kollektivavtalet.
Adressen är Mejlansvägen 2.
Som företagare till Finland:
Anvisningarna för sorteringen skiljer sig något från varandra i olika delar av landet.
Läs mer: Hobbyer för barn och unga
Löneanspråket får inte vara för stort, men inte heller för litet.
När du letar efter en hyresbostad kan du leta efter annonser till exempel på internet.
Personer som uppträder i videoklippet och tillstånd
Om du har ett körkort som utfärdats i ett land som inte är anslutet till Genève- eller Wien-konventionerna kan du köra bil med detta kort under ett års tid efter att ha registrerats i befolkningsregistret i Finland.
Finlands Konsumentförbunds rådgivningstjänst:
Ungdomsgårdar och -lokaler finska _ svenska
Tfn 044 977 4547
Mer information finns på Aalto-universitetets, Laureas och Metropolias webbplatser.
Uppgifterna om barnets födelse skickas från sjukhuset till befolkningsdataregistret i Finland.
Förälder eller annan vårdnadshavare
Finskundervisning ges på daghem, i förskola och skola.
Barn och motion
Information om social kreditgivningfinska _ svenska _ engelska
Invandrarelever använder i huvudsak grundskolans och gymnasieskolans vanliga tjänster.
Kurser hålls på finska, engelska och ryska.
Information om löneutbetalningfinska _ svenska _ engelska
I Helsingfors finns många simhallar, gym, idrottsplatser och motionsspår.
Hjälp med babyn
Då kan barnet även lära sig finska eller svenska som andra språk, som S2-språk (S2-kieli).
Kom ihåg att uppdatera din ansökan när den är i kraft. Annars löper den ut.
Läkaren bedömer din rörelsenedsättning och därefter kan du få hjälpmedel i form av medicinsk rehabilitering.
Läs mer på InfoFinlands sida Stöd- och serviceboende.
På internet finns många annonser om bostäder som är till salu.
Skatt betalas på alla arbetslöshetsförmåner.
Du hittar mer information på föreningens webbplats på finska, svenska och engelska.
I ett nytt företag uppskattar företagaren själv storleken av den beskattningsbara inkomsten och meddelar denna till skattmyndigheten.
Hiihtomajantie 2
Banken har även rätt att kontrollera om du har betalningsanmärkningar.
Om man inte har uppgjort ett skriftligt arbetsavtal ska arbetsgivaren utan särskild begäran ge en skriftlig redogörelse för de centrala villkoren i arbetet.
Privata tandvårdstjänster
Du kan inte få en finsk personförsäkring om du inte omfattas av den sociala tryggheten i Finland.
Du måste betala avgiften när du lämnar in ansökan om uppehållstillstånd.
På rådgivningsbyrån (neuvola) följs hälsa och uppväxt bland barn under skolåldern.
återflyttning
I den förberedande utbildningen läser barnen det finska språket och grundskolans läroämnen.
Om du har ett bibliotekskort kan du också använda internet gratis på biblioteken.
Skolor kan ha till exempel följande inriktningar:
Mer information om tjänsterna för handikappade hittar du på Esbo stads handikappservice.
Här finns böcker, musik, tidningar och tidskrifter samt ljudböcker på flera olika språk.
Gemensam ansökan till universitetfinska _ svenska
Om du behöver preventivmedel eller abort eller misstänker att du har en könssjukdom, kan du kontakta preventivmedels- och familjeplaneringsrådgivningen.
Esbo stad ordnar olika tjänster för handikappade, till exempel dagverksamhet och färdtjänster.
Hälsovården besöket barnet också hemma direkt efter födseln.
Till hemfrid.
Före äktenskapet ska du skriftligt begära hindersprövning (avioliiton esteiden tutkiminen).
När du ansöker om registrering av uppehållsrätt, kan du på samma blankett också begära att få en finsk personbeteckning.
Du kan ansöka om tjänster och stödfunktioner hos stadens socialarbetare.
De flesta tidningarna är finskspråkiga.
Om ditt boende i Finland inte anses stadigvarande, kan du ändå ha rätt att omfattas av den sociala tryggheten i Finland på grund av att du arbetar.
Fristående examina kan avläggas vid yrkesläroanstalter och vuxenläroanstalter.
Behovsprövad rehabilitering
hälsovård
Telefon: 040 193 6468
Läs mer på InfoFinlands sida Företagsrådgivning.
Några lagar
Rovaniemi regiontaxi erbjuder taxitjänster i Rovaniemiområdet dygnet runt.
Vi skickar ut korta webbenkäter högst varannan månad som rör innehållet i InfoFinland, webbplatsen eller kommunikation.
Om du äger en bostadsaktie betalar du vanligen
Du kan också bo som gäst hos vanliga finländare.
Fiske och båtlivfinska
bostadslånets storlek
Settlementföreningen Rovalan Setlementti ry/MoniNet
om du vill bli antagen för studier i ett visst ämne vid en högskola
På Grankulla stads webbplats kan du skicka respons till förvaltningen.
Mariegatan 28
I Helsingfors finns tre TE-byråer.
Du kan ansöka om registrering av uppehållsrätten om din försörjning i Finland är tryggad.
Familjen kan själv be barnskyddsmyndigheterna om hjälp.
Vad bör jag beakta innan jag undertecknar hyresavtalet?
Vad gör jag om det börjar brinna hemma?
Du kan göra en bostadsansökan på VAV Asunnot Oy:s webbplats.
Du måste även skaffa dig en bärbar dator.
Läs mer: Hälsa.
Esboområdet var bebott redan för ungefär 8 000 år sedan.
turism- och kosthållsbranschen
Enklast hittar du information om biograferna i ditt område, bioprogrammet och biljettpriserna på internet.
Dessa tjänster inkluderar bland annat:
Karleby huvudhälsostation
Du måste begära ett europeiskt recept särskilt av din läkare.
registreringsintyget över uppehållsrätten (om du är EU-medborgare)
Din skolresa måste vara minst 10 kilometer lång och resekostnaderna måste överstiga 54 euro per månad.
Om du inte behöver brådskande vård kan du tvingas vänta flera månader på en tid.
Man kan också flyga till många städer.
Anonyma narkomaner
Om du kommer till Finland för att arbeta under fyra månader, kan du ha rätt till hemvårdsstöd för barn och den offentliga hälsovården.
Nybörjarkurs i finska, Uunofinska
Esbo social- och krisjour
Om du är medborgare i ett nordiskt land och flyttar till Finland ska du registrera dig vid magistraten.
Upphovsmannen/den ansvariga personen ansvarar för alla eventuella upphovsrätts- och lagringsavgifter och rättsliga krav från tredje parter.
linkkiArbetslöshetskassornas samorganisation:
När du tar hand om en anhörig i hemmet
Läs mer på InfoFinlands sida Jämlikhet och jämställdhet i arbetslivet.
Arbetstagaren och den sociala tryggheten i Finlandfinska _ svenska _ engelska
Hur sopsorterar jag rätt?
Till exempel FPA (Kela) och Migrationsverket (Maahanmuuttovirasto) bokar i vissa situationer en tolk för klienten.
Om du flyttar till Finland för att bo här stadigvarande i minst ett år ska du också registrera dig som invånare i magistraten.
Du kan studera vid öppna högskolor
Om du till exempel har ett företag som idkar skönhetsvård eller säljer livsmedel ska företagets lokaler kontrolleras.
När du ringer nödnumret 112:
I kollektivtrafikens färdmedel kan du betala med kontanter eller resekort (matkakortti).
Läs mer om upprättandet av arbetsavtalet på InfoFinlands sida Innehållet i arbetsavtalet.
Arbetsgivarna ordnar utbildning i första hjälpen på arbetsplatsen.
Äktenskapslagenfinska _ svenska _ engelska
Fråga din chef hur långa pauser du har.
När du ansöker om finansiering måste du ha en ordentlig affärsverksamhetsplan färdig.
Fråga närmare uppgifter om undervisningen vid närmaste sommaruniversitet.
Om du känner att du inte klarar dig med babyn utan hjälp kan du bo på ett mödrahem och lära dig hur du tar hand om barnet där.
Järnvägsstationen finns i stadens centrum.
Navigatorn ger dig råd om utbildning, arbete, vardagen och livet.
Hotellfinska _ svenska _ engelska _ ryska
Familia Clubs projekt Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska.
Om äktenskapet slutar med att en av makarna dör, delas makarnas sammanlagda egendom mellan arvingarna till den avlidna makan och den maka som fortfarande lever.
linkkiAFAES:
Rätt att arbetafinska _ svenska _ engelska
Till de öppna högskolorna ordnas inga inträdesprov.
Finlands beskickningar utomlands
upphör när grundskolans lärokurs har fullgjorts eller det har förflutit 10 år sedan läroplikten började.
I Vanda finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
I Finland måste bilen besiktigas och registreras.
På rådgivningen följer man med moderns, barnets och hela familjens välmående under graviditeten.
Röda Korset ger också rådgivning om reglerna för familjeåterförening och därom, hur familjemedlemmarna ska gå tillväga för att ansöka om familjeåterförening.
Om du vistas i Finland tre månader utan avbrott behöver du inte ansöka om registrering av uppehållsrätten.
Läs mer: Motion.
Invandrare och grundläggande utbildning
Haartmansgatan 4
Samtala på finska
I höghus finns ett nummer nära entrédörren som du kan ringa i en sådan situation.
Språkstudier som arbetskraftsutbildning
Då behöver du inte heller betala mäklararvode (välityspalkkio).
Du hittar bostäder som hyrs ut av företag och privatpersoner via bostadssidor på internet.
linkkiMannerheims barnskyddsförbund:
linkkiApotekareförbundet:
Om uppehållstillståndet beviljats på någon annan grund än internationellt skydd, kan andra anhöriga inte få uppehållstillstånd.
Kontrollera att frånluftsventilerna är öppna.
familjens storlek och
Läs mer på InfoFinlands sida Barnbidrag.
Det finns ingen särskild asylansökningsblankett som du skulle kunna fylla i förväg.
I en del situationer kan myndigheten beställa en tolk och betala för tolkningen. Detta är inte alltid möjligt.
I Helsingfors finns det också många privata tandläkare.
När du flyttar utomlands måste du meddela detta till FPA, om du får FPA:s förmåner eller om du har det europeiska sjukvårdskortet.
På trafikverkets webbplats finns kollektivtrafikens reseplanerare, matka.fi, där du kan söka den bästa rutten och det bästa resesättet.
För att kunna göra det behöver arbetsgivaren ett skattekort av dig.
Kontaktuppgifter till skyddshemfinska _ svenska
integrationsutbildning
Ta med dig identitetsbevis och ett foto när du ansöker om kortet.
linkkiVasa ortodoxa församling:
Den evangelisk-lutherska kyrkan har fyra finskspråkiga församlingar och en svenskspråkig församling i Karleby.
På många jobbsajter kan du spara din jobbansökan och meritförteckning (CV) så att arbetsgivaren kan läsa dem.
Flera av Matkahuoltos bussar i lokal- och regiontrafiken avgår från Rovaniemi busstation.
Har du rätt till förmåner?
Om det inte hjälper, kontakta arbetsplatsens förtroendeman.
Finlands Konsumentförbund erbjuder råd och handledning både för hyresgäster och hyresvärder.
Båtlivfinska _ svenska _ engelska
Den katolska kyrkan kom till Finland via Sverige och den ortodoxa kyrkan från Novgorod i öster, nuvarande Rysslands område.
Utbildningsavtalet kan även kombineras med läroavtal.
Det finns också andra villkor; till exempel måste du kunna visa hur du försörjer dig.
_ litauiska
I Finland föder de flesta mammor vaginalt.
Till exempel ska man ha varit med i arbetslöshetskassan en viss tid före man blir arbetslös.
Arbetsgivaren är skyldig att teckna pensionsförsäkring åt alla sina anställda och betala försäkringspremierna.
Steinergymnasietfinska
Finland under vistelsen och inte stannar i landet tre månader utan avbrott, behöver du inte ansöka om registrering av uppehållsrätten.
Helsingfors-Vanda internationella flygplats ligger i Vanda.
Finland har ingått avtal om den sociala tryggheten med ett antal länder.
Information om Helsingfors(pdf, 5,9 MB)finska _ svenska _ engelska _ ryska _ franska _ kinesiska _ tyska
Familjerådgivningar och familjecenter finns på många orter.
Stöd kan betalas till en person eller till ett hushåll (ruokakunta).
Hälsostationerna enligt stadsdelfinska _ svenska _ engelska
Vänligen observera att endast Migrationsverket kan fatta beslut om uppehållstillstånd.
Vid Grankulla medborgarinstitut kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Rådgivning för invandrarefinska
Arbetspensionsförsäkringsbolag, pensionskassor och -stiftelser har hand om arbetspensionsförsäkringarna.
Intressebevakning och rådgivning för företagare
yrkeshögskolan Laurea
Som företagare betraktas:
Rabatt på bussbiljetter ges åt
Under kvällar och helger är hälsostationerna stängda.
Stöden för pensionärerfinska _ svenska _ engelska
Sommaruniversitetet
När ansökan avgjorts, ser du beloppet på ditt stöd och tidpunkten för utbetalningen.
Den sociala tryggheten
I Grankulla anordnas förskoleundervisningen i daghemmen.
Innan du kan få ett uppehållstillstånd måste du hitta ett jobb i Finland.
Den evangelisk-lutherska och den ortodoxa kyrkan har en särställning i Finland.
Information och hjälp för rusmedelsberoendefinska _ svenska _ engelska _ ryska
Den är avsedd för stadens invånare.
Hälsostationernas kontaktuppgifter finns på Esbo stads webbplats.
Seniori-info
Den avlidne kan ibland ha rätt till begravningsbidrag (hautausavustus) genom sitt senaste anställningsförhållande eller medlemskap i ett fackförbund.
Du ska alltid först ansöka om grundläggande utkomststöd hos FPA.
Skolan börjar (läroplikt).
linkkiEsbo musikinstitut:
Utöver stadens egna skolor finns det privata skolor och statliga skolor i Helsingfors.
Hemvårdsstöd
En delägarbostad (osaomistusasunto) är ett bra sätt att skaffa en egen bostad om du inte kan köpa dig en egen bostad direkt.
Gymnasium och yrkesläroanstalt
Information om tandvården för skolbarnfinska
1812 Helsingfors blir huvudstad
Moderskapsförpackningen innehåller bebiskläder och vårdartiklar.
Det är relativt dyrt att köpa och använda en bil i Finland.
Då utför du praktiska arbetsuppgifter i verkliga situationer på en arbetsplats.
Du får även stöd när du funderar på om du ska starta ett företag.
Information om stadenfinska _ svenska _ engelska
I Finland utgår man alltså inte från att enskilda människor tar hand om sådana släktingar som har det dåligt ställt ekonomiskt.
Om barnet inte får finskt medborgarskap
Undervisningsspråket i vid Karleby finska gymnasium och Karleby vuxengymnasium är finska och svenska vid Karleby svenska gymnasium.
inte uppfyller villkoren för inkomstrelaterad dagpenning.
Grunderna för FPA:s bidrag definieras i lagen.
År 1995 blev Finland medlem i Europeiska unionen (EU).
Språkexamen finns på tre olika nivåer: för nöjaktiga, goda och utmärkta språkkunskaper.
Stöd för vård av en handikappad anhörig
Beloppet på din föräldradagpenning beror på hur höga inkomster du har.
Vid skilsmässa eller när sambor flyttar isär måste föräldrarna besluta om barnets vårdnad, underhåll, boende och umgängesrätt.
Magistraten i Nyland, Esbo enhet
Om du behöver hjälp eller råd i skötseln av dina personliga ärenden, ta då direkt kontakt med myndigheterna.
Om du har en utländsk examen
Kulturevenemang för barnfinska
Abiturientkurser (abikurssi) för gymnasieelever som förbereder sig för studentskrivningarna
Socialhandledare 016-322 3125, 040-576 8904
Läs mer på InfoFinlands sida Integration i Finland.
I Finland är våld brottsligt.
anställningsform
Jouren är avsedd för patienter vars sjukdom kräver brådskande bedömning och vård.
Finland finansierade tillverkningen av varorna med lån och understöd.
Många bor också långt från centrum eller i en närliggande kommun och pendlar långt till jobbet.
Flera olika föreningar samt kommunala institut ger unga möjlighet att studera idrott och kultur samt bl.a. språk och hantverk.
Lapplands arbets- och näringsbyrå
Högst är priserna i centralt belägna bostäder.
Specialvårdspenning för barn under 16 årfinska _ svenska _ engelska
Vad är ditt telefonnummer / din e-postadress?
Barnatillsyningsmannen
Du måste studera på heltid.
Mer information hittar du via tjänsten Helsingforsregionen.fi.
Tidningar
Det är också viktigt att känna till sina kunder och försäljningsmetoder.
Information om högre yrkeshögskoleexamenfinska _ svenska
FPA sköter folkpensionerna och garantipensionerna.
Skatteprocenten på kapitalinkomsten är alltid densamma.
Mer information hittar du på organisationens webbplats.
Arbetslivet i Finland styrs av många regler som arbetstagaren och arbetsgivaren måste följa.
Simning och skidåkning är mycket populära grenar i Finland och i dem ordnas nybörjarkurser även för vuxna.
Lapplands regionkontor/ Rovaniemi serviceställe
Barnskyddet är baserat på barnskyddslagen och internationella konventioner.
Skriv ett eget CV för varje arbetsplats.
Information om Finlands Dövas Förbundfinska _ svenska _ engelska
Mottagningspenningen är ett litet belopp som är avsett för ofrånkomliga utgifter.
I Karleby finns hälsostationer i olika delar av staden.
Om du behöver brådskande hjälp av polisen, ring nödnumret 112.
Din uppehållsrätt kan registreras om du har en familjemedlem som är stadigvarande bosatt i Finland.
Läs mer: Småbarnspedagogik
Strandgatan 16 (våning 5 och 6)
Hyresbostäder för studerande erbjuds av Helsingforsregionens studentbostadsstiftelse HOAS och Aalto-universitets studentkår AUS.
Telefontid och tidsbokning
Öppningsoperationen kan även göras i mitten av eller före graviditeten.
Dessutom utreder ditt ombud om du kan återförenas med din familj.
Rättighet:
I Rovala-institutets utbildning för invandrare kan man studera det finska språket och den finska kulturen, arbetslivsfärdigheter och skaffa sig kunskaper om det finländska samhället.
Studierna är allmänbildande: fokus ligger speciellt på naturvetenskapliga och humanistiska ämnen.
Om du är ung kan du berätta om det som bekymrar dig till exempel för skolhälsovårdaren, skolpsykologen eller skolkuratorn.
Vigselfinska _ svenska _ engelska
Faderskapet kan fastställas vid mödravården under graviditeten.
kan fadern vara barnets vårdnadshavare antingen tillsammans med barnets mor eller ensam.
Logga in med nätbankskoder eller ett mobilcertifikat.
Till gymnasieutbildning för ungdomar ansöker man under våren via gemensam ansökning för gymnasierna och man kan bli antagen om man i slutbetyget från grundskolan har tillräckligt högt snittbetyg i läsämnena.
Öppettider: mån-fre 9-17
Socialbyrån
Grundundervisning för vuxnafinska
Information om busstidtabellerna hittar du på Matkahuoltos webbplats och verksamhetsställen.
Medelnivån är avsedd för personer som kan språket relativt väl. Deras färdighetsnivå är 3–4.
Enligt lag ska arbetsgivaren betala högre lön för övertid.
Familjebandet mellan föräldern och barnet måste bevisas, till exempel med en födelseattest med föräldrarnas namn.
Prövningen görs vid magistraten. Du kan lämna in ansökan om prövning vid vilken magistrat som helst.
Annan anhörig till en finsk medborgarefinska _ svenska _ engelska
Läs mer: Problem i äktenskap och parförhållande
Ibland behövs det skrapning efter medicinsk abort.
Hyresnivån är hög i Helsingfors.
Dessutom krävs det att familjelivet upphört på grund av ett tvingande skäl, till exempel för att man blivit flyktingar.
Besöksadress: Karlebygatan 27, Karleby
Se till att du har försäkringar.
I vissa fall får du tolken via myndigheten.
De flesta arbetsgivare värdesätter att den anställda vill utveckla sig i sitt arbete och inhämta nya kunskaper.
Inte heller intyg som utfärdats av en ambassad eller ett konsulat i Finland behöver legaliseras.
År 1920 blev villasamhället en köping.
Skilsmässa utan betänketid
Om du lider av en yrkessjukdom eller har blivit skadad i ett olycksfall, kan du få rehabilitering från försäkringsbolaget (vakuutusyhtiö).
linkkiVästra Nylands rättshjälpsbyrå:
Nuppi
I sådana situationer avvägs alltid fall till fall om uppehållstillståndet förlängs efter skilsmässan eller om det återkallas.
Du kan ringa jourtelefonen dygnet runt.
Strandgatan16
Information om den sociala tryggheten i Finlandfinska _ svenska _ engelska
Film, dans och teaterfinska _ engelska
Vanda stad betalar dessutom ett kommuntillägg till hemvårdsstödet för barn till de familjer som vårdar ett under 1 ½-årigt barn i hemmet.
Familjerådgivningscentralen vid Rovaniemi församling
Läs mer: Motion.
ogifta barn under 18 och deras vårdnadshavare som bor i Finland
Finlands Näringsliv EK representerar alla privata branscher och företag i alla storlekar.
Lediga tjänsterfinska
Alla som ansöker om en förskoleplats ska lämna in en ansökan om förskoleundervisning.
I vissa fall behövs det dock ett tillstånd från myndigheter för att starta företagsverksamhet, eller också måste man anmäla verksamheten till myndigheter.
Fristående examen (näyttötutkinto) är ett sätt att bevisa sin yrkeskunnighet.
Arbetskraftsutbildning är i huvudsak utbildning avsedd för arbetslösa arbetssökande.
I Helsingfors finns många olika religionssamfunds tempel och dessutom olika verksamhetscenter.
Du kan få full arbetslöshetsförmån om du under 65 betalningsdagar, alltså under cirka tre månaders tid, utför en viss mängd lönearbete, får inkomst som företagare eller deltar i en verksamhet eller en tjänst som främjar din sysselsättning.
linkkiKärlek och anarki:
Gå igenom dina utbildningar och din arbetserfarenhet och fundera på vilka färdigheter du lärt dig i dem.
Utkomstförutsättningfinska _ svenska _ engelska
Du behöver en personbeteckning när du sköter ärenden hos myndigheter, och dessutom underlättar den skötandet av ärenden i till exempel banker och med din arbetsgivare.
På InfoFinlands sida Familjemedlem finns mer information för dem som flyttar till Finland på grund av familjeskäl.
När du har fått ett positivt utlåtande från Business Finland kan du ansöka om uppehållstillstånd för uppstartsföretagare hos Migrationsverket.
Yrkesläroanstalterfinska _ engelska
Byrån i Esbo finns i Alberga.
Statens lokalförvaltningfinska _ svenska
Prövotid och längden på den
Från och med den 1 april 2019 kan studerande från länder utanför EU och EES ha rätt till vissa förmåner, till exempel förmåner som ingår i sjukförsäkringen.
Läs mera på InfoFinlands sida Bostadsbidrag.
Ett nödfall är en verklig och akut farlig situation där ens liv, hälsa, egendom eller miljön är hotad.
Barnets sociala trygghet
Hen hjälper elever som har det svårt i skolan.
Per telefon betjänar socialjouren och krisjouren på finska, svenska och i mån av möjlighet även på engelska.
Vi följer automatiskt besökarna i tjänsten och använder informationen till att utveckla tjänsten.
Teckna en pensionsförsäkring senast när det har gått sex månader sedan du startade företagsverksamheten.
Arbete och entreprenörskap
Ansökningsblanketterna kan hämtas från och lämnas in till Kokkolan Vuokra Asunnot Oy:s verksamhetsställen.
Barnförhöjningfinska _ svenska _ engelska
Barn, vars föräldrar har skilt sig, har rätt att vägra träffa någon av föräldrarna.
För att få inkomstrelaterad dagpenning finns några villkor som måste uppfyllas innan det är möjligt att få dagpenning.
När man har avlagt magisterexamen, kan man ansöka om rätt till fortsatta studier och avlägga licentiat- eller doktorsexamen.
Undervisning för invandrare
linkkiTukes:
Information om öppna universitetetfinska _ svenska
Telefonen betjänar på finska, svenska, engelska och tyska.
Pass
du är av finländsk härkomst
Tfn 040 701 8446
I utrustningen i en hyresbostad ingår nästan alltid köksskåpen, kylskåpet och spisen.
Stadens borgare köpte tjära av bönder och exporterade den, ofta till hamnar vid Medelhavet och i England.
Webbplats för Asokoditfinska
Helsingfors ungdomsstation (Helsingin nuorisoasema) erbjuder hjälp till 13–23-åriga unga Helsingforsbor.
I förskolan lär sig barnen att uppskatta sitt språk och sin kultur.
Sådan verksamhet ordnas till exempel av församlingar och organisationer.
Att grunda ett företag
Stöd för unga invandrarefinska
Sökning av relationsrådgivningstjänsterfinska _ svenska _ engelska
I de större parkerna kan man övernatta och göra längre utflykter.
Du kan be om råd per telefon (06) 826 4477.
Senare blev Kokkola stadens finska namn.
Museisökningfinska _ svenska _ engelska
fre kl. 8–14
Stadens hyresbostäder
linkkiFöretagarna i Finland:
Om du blir kallad till hälsovården, kom ihåg att på förhand ange att du behöver en tolk.
Parförhållande
linkkiSHVS:
Hyresbostäder för personer under 30 årfinska _ engelska
Med ett rasistiskt brott avses ett brott som förövaren begår av rasistiska orsaker.
Utbytesstudenter
Studiebostäder hyrs ut av Kiinteistöyhtiö Tankkari, som erbjuder möblerade kollektivbostäder samt familjebostäder i olika storlek.
Kontakta ditt försäkringsbolag direkt när skadan har inträffat.
Karleby evangelisk-lutherska församlings arbete bland missbrukarefinska _ svenska
Grankullavägen 10
Utbildning i finska och svenska språketfinska _ svenska _ engelska
När du tar emot en studieplats, förbinder du dig att börja studera i läroanstalten.
De berättar inte om dina saker för andra myndigheter.
Grankullas areal är 6,0 km2.
En del teatrar är professionella, andra är amatörteatrar.
1523 Gustav Vasa blev kung över Sverige och lösgjorde Sverige från den medeltida nordiska unionen.
Du får ett nytt skattekort:
Företagandet kan också upphöra om företaget säljs, avvecklas, går i konkurs, försätts i likvidation eller på grund av skilsmässa.
Stöd för närståendevårdfinska
Vanligen är hyrestiden ca 5-12 år.
På stadens webbplats hittar du också anvisningar om hur du söker hyresbostad.
Finlands Rösa Kors hjälper med researrangemangen för kvotflyktingar
bor stadigvarande i Finland
Biobiljetternas priser varierar något i Finland.
Kultur för barn och ungafinska _ svenska _ engelska
Flytt utomlands och den sociala tryggheten
Orsaken till barnlöshet kan finnas hos kvinnan eller hos mannen.
Ansökan kan lämnas till tingsrättens kansli eller skickas dit per post, fax eller via e-post.
Identitetskort för utlänningar
När hyresgästerna väljs beaktas
Adress: Östersjögatan 3
Också föreningar och idrottsklubbar ordnar mycket verksamhet för ungdomar.
Du hittar kontaktuppgifterna på Håkansböle internationella förenings webbplats.
Uppehållskort för en familjemedlem till en EU-medborgare
Tfn (09) 8392 4342
Om barnet flyttar till Karleby under läsåret kan han eller hon genast börja i skolan.
Du kan söka folkpension och garantipension om du omfattas av Finländska socialskyddet och när du har bott i Finland minst tre år efter att du fyllde 16 år.
Arbetarskyddsmyndigheter
Som ensamstående förälder har man själv ansvaret för fostran av barnet.
linkkiFöreningen för familjer med en förälder r.f.:
arbetspraktik som ingår i examen eller ett slutarbete eller
Du kan boka en tid på Migrationsverkets tidsbokningstjänst.
Om du bor i Helsingforsregionen, Tammerforsregionen eller Åboregionen kan du leta efter en kurs i finska språket som passar dig genom tjänsten Finnishcourses.fi.
Hälsostationen på Pulkamontiefinska
Det finns två slags resekort.
Pensionsförsäkringen tryggar företagarens utkomst då företagsverksamheten upphör på grund av invaliditet eller ålder och den ger företagarens anhöriga ett familjepensionsskydd efter att företagaren har dött.
Om du har kraftiga smärtor eller blödningar ska du kontakta sjukhuset.
Du kan ansöka från Kela om ekonomiskt stöd för hemvård av barn.
Om du vårdar ditt barn hemma även efter detta har du rätt att vara ledig från ditt arbete för vård av barn tills barnet fyller tre år.
Idrottsanläggningar
linkkiDidar:
Om barnet inte har tillräckligt bra kunskaper för att klara grundskolan kan han eller hon få förberedande undervisning.
Realämnen (reaali), d.v.s. historia, religion, fysik, kemi, biologi, psykologi, filosofi
Om du själv bokar tolken och betalar kostnaderna, kan du anlita en tolk när som helst.
När barnet fyller två år kan du inte längre ta ut faderskapsledighet trots att du har dagar kvar.
I Finlands finns ungefär ett tusen museer, varav cirka 300 är regelbundet öppna för allmänheten.
Du kan ansöka om tillståndet elektroniskt via tjänsten Enter Finland eller på Migrationsverkets tjänsteställe.
Mödrarådgivningen ger alla blivande föräldrar broschyren Vi väntar barn som ges ut av Institutet för hälsa och välfärd (Terveyden ja hyvinvoinnin laitos).
Info om HIVfinska _ engelska _ ryska
Fordon som flyttgodsfinska _ svenska _ engelska _ ryska
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åriga ungdomar.
Pyrolavägen 37
Information om barnskyddfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Integrationen underlättas t.ex. av att
linkkiÖstra Nylands rättshjälpsbyrå:
Om du inte kan något av dessa språk, ska du fråga om det är möjligt att anlita tolk när du bokar tid till tandvården.
linkkiFFC:
Kriscentret vid Lapplands mödra- och skyddshem
Invandrare som har bott tillräckligt länge i Finland får ålders- eller invalidpension på samma grunder som alla andra som är bosatta i Finland.
Ruttkartor säljs i bokhandlar och på internet.
Studier i finska språket på Internetfinska _ engelska
Om du är över 65 år kan du kontakta seniorrådgivningen vid Grankulla hälsostation.
Svenska är modersmålet för cirka 5 procent av finländarna.
Vanligen motsvarar garantin beloppet på två månaders hyra.
Planeringen och konstruktionen av kärnkraftverket är ett omfattande projekt som tar cirka 10 år att slutföra.
Du kan tillförlitligt intyga din identitet.
Stödcentret betjänar alla, oavsett kön.
Du kan också söka skilsmässa ensam, utan din makes eller makas samtycke.
Festivalerna ordnas på olika håll i Finland, både i städerna och på landsbygden.
För detta behövs dock ett undervisningstillstånd från Trafi.
Barn med invandrarbakgrund kan få undervisning i det egna modersmålet.
Vid Lapplands yrkesinstitut kan du studera och skaffa dig yrkesinriktad grundutbildning och vuxenutbildning i alla studieområden förutom inom idrottsområdet och turism-, kosthålls- och ekonomibranschen.
Information om hur du ansöker om tillståndet finns under rubriken Att ansöka om uppehållstillstånd.
I Finland finns det 24 flygplatser.
Förskoleundervisning
Du kan få fortbildning eller påbyggnadsutbildning i din egen bransch.
Till följd av Sovjetunionens kollaps och den ekonomiska tillväxten på 1980-talet som baserade sig på lån hamnade Finland i depression på 1990-talet.
Mer information om anmälan får du på Utbildningsstyrelsens (Opetushallitus) webbplats.
Kontaktuppgifter
Information om utkomststödfinska _ svenska _ engelska
Försörjningsförutsättningen gäller er även i det fall att ni gifte er efter att din make/maka kom till Finland.
om du tar hand om barnet i hemmet och hemvården ansluter sig till barnets sjukhusvård eller
Ett brottmål kan även medlas, om offret och den brottsmisstänkta samtycker till detta.
Under kvällar och veckoslut finns tandvårdsjouren (hammashoidon päivystys) vid Haartmanska sjukhuset i Helsingfors.
Också parets gemensamma barn kan bo med familjen.
Föreningen för bostadslösafinska
Studentkåren vid Lapplands universitet informerar också om bostäder som hyrs ut till studerande.
Trafiken i Finland.
Fråga mer av läkaren vid din egen hälsostation (terveysasema).
De vill dessutom stärka InfoFinlands riksomfattande ställning, så att det är möjligt för nya kommuner och andra organisationer att ansluta sig till tjänsten också i fortsättningen.
Att bli av med sin bostad
Efter betänketiden
Dessutom är det även möjligt att läsa normala gymnasiekurser vid sommaruniversitetets sommargymnasium.
När du går till TE-byrån ska du ta med dig
Beslutsfattandefinska _ svenska _ engelska
Upphovsmannen som deltar i tävlingen överlåter till tävlingsarrangören, Helsingfors stad, obegränsad rätt att kostnadsfritt visa verket offentligt och att utnyttja verket eller delar av verket i sin marknadsföring av Infobanken på Internet och i andra motsvarande medier samt internationella evenemang.
Information om företagarpensionsförsäkringenfinska _ svenska _ engelska
Hjälp till offer för människohandelfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ thai _ vietnamesiska _ polska _ rumänska _ bulgariska
Dessutom erbjuds åldringar i Esbo egna tjänster, till exempel hemvårdens tjänster.
Bostaden kan till exempel byggas om så att du kan röra dig med en rullstol i den.
Du betalar samma skatt hos alla dina arbetsgivare.
Den avlidne kan begravas i kista eller kremeras.
Musikundervisning för barn och vuxnafinska _ engelska
Antalet kommunfullmäktige beror på kommunens invånarantal.
Yrkesinriktad grundexamen
linkkiYle:
Typiska ledda aktiviteter är olika temadagar och utflykter.
På biblioteket kan du låna böcker på klarspråk som är skrivna på lättläst finska.
Skilsmässa i ett bikulturellt äktenskapengelska
Utbildning som handleder för grundläggande yrkesutbildning (Ammatilliseen peruskoulutukseen valmentava koulutus) d.v.s. VALMA är avsedd för dem som vill avlägga en grundläggande yrkesutbildning.
Om du skiljer dig på grund av att din make/maka varit våldsam mot dig kan ditt uppehållstillstånd förlängas trots skilsmässan.
Du kan få startpenning för högst tolv månader.
Elarbeten som du får göra självfinska
Om du ansöker om fortsatt uppehållstillstånd först efter att ditt tidigare uppehållstillstånd gått ut, får du uppehålla dig i Finland under tiden då ansökan behandlas men har inte rätt att arbeta innan du erhållit fortsatt uppehållstillstånd.
Tfn 09-228 05141, mobil 050 325 7173 (ryska, engelska)
Du ingår ett avtal med företaget och företaget skickar dig till arbete för en annan arbetsgivare.
ons–fre kl. 17–21
Du ansöker om visum i den närmast belägna finländska beskickningen eller visumcentralen.
Alla texter som publicerats på InfoFinlands webbplats på alla språk är fritt tillgängliga i enlighet med licensen Creative Commons Erkännande 4.0.
Om du är frånskild kan du gifta om dig utan tillstånd från din före detta maka eller make.
Serviceboende
integrationstjänster
Fågelbergavägen 2 A
Hjälpmedel kan fås tidigast när barnet går i grundskolans årskurs sju.
Skilsmässa i Finlandengelska _ ryska _ estniska
Du kan ringa A-klinikens medarbetare mån–fre kl. 8.30–10, tfn 040 195 3981
Många företag gick i konkurs, vilket fick till följd att många människor förlorade sina jobb.
Om du behöver mer krävande vårdåtgärder, som till exempel tandkirurgi, ska du först boka tid hos en tandläkare.
Du kan ansöka om utbetalning av arbetslöshetsersättning till Finland med blankett E303 eller U2.
Det finns även många organisationer där du kan få information och stöd.
du har anmält dig som arbetssökande vid arbets- och näringsbyrån och din jobbsökning är i kraft
Arbetslivets ABC finska
Utbetalning av pension till utlandet
Information om FPA:s hemvårdsstödfinska _ svenska _ engelska
Du behöver ingen remiss till A-kliniken, utan kan själv boka en tid.
Regeringen (hallitus) består av statsministern och de andra ministrarna.
Kom i tid till mottagningen.
Fråga den senaste arbetsgivaren eller fackförbundet om detta.
I Helsingfors finns även många invandrarföreningar.
Du kan använda tjänsten på finska, engelska och ryska.
Tjänsten är finskspråkig.
Släng inte föråldrade läkemedel utan lämna dem alltid till apoteket (apteekki), eftersom de är problemavfall.
Tack vare det effektiva biblioteksnätverket i Finland är nästan alla finländska biblioteks samlingar tillgängliga för bibliotekskunderna i Karleby.
Det är bra att upprätta ett skriftligt avtal om underhållsbidraget som socialnämnden bekräftar.
Domstolen dömer till skilsmässa först efter att den andra ansökan har lämnats in.
Arbeta i Finland
Du kan söka till många olika läroanstalter i den gemensamma ansökan.
Medborgare i EU-länderna, Island, Liechtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns nättjänst.
Boendeservice för utvecklingsstördafinska
Duo erbjuder relationsrådgivning för par från två kulturer på finska och engelska.
Tidpunkten då arbetet inletts
Denna lag tillämpas bland annat på diskriminering på grund av etniskt ursprung inom offentliga och privata social- och hälsovårdstjänster.
Kollektiv- och tjänstekollektivavtalet är bindande för de löntagar- och arbetsgivarförbund som slutit dem och för deras medlemmar.
Förskoleundervisning (esiopetus) ordnas i både kommunala och privata daghem samt i förskoleenheter i skolornas lokaler.
Omskärelse av kvinnor och flickorfinska _ engelska _ somaliska _ arabiska
Anmäl flyttningen till myndigheterna
Integration av och rådgivning för invandrare
Mer information om medling i familjefrågor får du på justitieministeriets webbplats.
I brådskande fall behöver du ingen remiss.
Om du misstänker att en arbetsgivare, en läroanstalt eller någon annan instans har diskriminerat dig på grund av ditt kön och brutit mot lagen om jämställdhet mellan kvinnor och män, kan du be jämställdhetsombudsmannen om råd och anvisningar samt hjälp med att utreda ärendet.
Lämna in din ansökan på internet i tjänsten Enter Finland eller vid Migrationsverkets tjänsteställe.
registrering av uppehållsrätten om du är EU-medborgare
När du går till magistraten ska du ta med dig åtminstone följande handlingar:
Du kan behöva intyget också när du söker ett jobb eller en studieplats.
Om du behöver rådgivning och handledning om integration kan du kontakta Rovaniemi stads integrationsrelaterade socialtjänster.
Om du behöver hjälp med att använda Wilma ska du be skolan om en introduktion.
du har ett tillfälligt uppehållstillstånd på grund av hinder för avlägsnande ur landet
Du får stanna i Finland om du beviljas asyl eller uppehållstillstånd på andra grunder.
Detta beror på huruvida det andra landet godkänner flerfaldigt medborgarskap för barnet.
maskiner och utrustning
kopia på uppehållstillstånd eller pass om du inte är EU-medborgare.
När barnet börjar i dagvården fyller man tillsammans med familjen i blanketten Uppgifter om invandrarbarn.
Även arbetsgivaren kan förutsätta att arbetstagaren inte har betalningsanmärkningar.
Skriv in sökordet ”hyresbostad”.
Håkansböle hälsostation, Galoppbrinken 4
Via tjänsten Uskonnot Suomessa kan du söka information efter det religiösa samfundet och orten.
Konserter ordnas på olika platser: I konsertsalar, musikhus, kulturcenter, institut, restauranger, på historiska platser och i kyrkor.
Uppehållskortet för en familjemedlem till en EU-medborgare beviljas för fem år eller en kortare tid om boendet i Finland varar mindre än fem år.
Medarbetaren vid servicestället kan hjälpa dig att fylla i ansökningen.
Den länsbaserade handredskapsavgiften är personlig och ska betalas innan fisket påbörjas.
Vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto) kan 17–24-åriga invandrarungdomar avlägga grundskolans avgångsbetyg.
Dessa länder är de nordiska länderna (Sverige, Danmark, Norge och Island), USA, Kanada och Quebec, Chile, Israel, Indien och Australien.
Kommunal småbarnspedagogik
Skolhälsovårdaren tar hand om skolbarns hälsa.
Du kan få hjälp med att överklaga av antingen en privat jurist, en statlig rättshjälpsbyrå (valtion oikeusaputoimisto) eller Flyktingrådgivningen rf (Pakolaisneuvonta) (endast asylsökande).
Arbets- och näringsbyråerfinska _ svenska
Du blir också tvungen att betala försäkringspremier, om du inte är försäkrad i det land där du bor stadigvarande.
Tillståndet kan beviljas om:
hur semestern bestäms
försäkringar
Du kan ansluta dig till ett fackförbund genom att ta kontakt med förtroendemannen på din egen arbetsplats eller genom att kontakta fackförbundet direkt.
Omskärelse av pojkar
Hotellfinska _ svenska _ engelska _ ryska _ kinesiska
tis–fre kl. 9–16, besök hos handläggarna endast med tidsbeställning
Examen är avgiftsbelagd.
Valmansföreningen ska ha minst 2 000 medlemmar.
För att få uppehållstillstånd på grund av familjeband måste du vara barnets vårdnadshavare.
Bostadsbidrag beviljas endast för skäliga boendekostnader.
Skatteförvaltningen räknar ut en lämplig skatteprocent åt dig utgående från hur mycket du förtjänade året innan.
har varit medlem i arbetslöshetskassan i minst 26 veckor innan du blev arbetslös.
Våld kan vara till exempel
Tfn 016 322 4900.
Läroplikten
Läs mer: Att röra sig i naturen.
Enligt lagen har barnets föräldrar eller vårdnadshavare huvudansvaret för barnets välfärd och harmoniska utveckling.
Tolktjänsterfinska _ svenska _ engelska
Studierna ska leda till
Om din make/maka/sambo/partner har fått flyktingstatus den 1 juli 2016 eller efter detta ska ansökan om uppehållstillstånd lämnas in inom tre månader efter att hen fått beslut på sin ansökan.
Allmänna språkexaminafinska _ svenska _ engelska
Hos Takuusäätiö kan du få hjälp och råd med betalningen av skulder.
Köp och konsumentens rättigheter
Språkexamen finns på tre olika nivåer: grundnivån, mellannivån och högsta nivån.
Snön smälter vanligen i mars eller april.
Läs mer: Föreningar.
På vissa arbetsplatser, till exempel sjukhus, arbetar man även under helgerna.
Information om sommaruniversitetetfinska _ svenska _ engelska
Vid val av invånare till stadens hyresbostäder prioriteras de sökande som har ett akut bostadsbehov.
Du ska också ha en arbetsplats som uppfyller kraven.
När du har en bostad är det bra att också ta en hemförsäkring (kotivakuutus).
För att få uppehållstillstånd för företagare måste du själv arbeta i ditt företag i Finland.
I Finland kan hälsovårdare ge vård vid flera sjukdomar.
Könssjukdomar behandlas på hälsostationen och på polikliniken för könssjukdomar i Helsingfors. .
Ansökan om hyresbostad i stadenfinska _ engelska
Skapa nätverk och upprätthåll ditt kunnande
Familjer kan få olika slags understöd för sina levnadskostnader.
Arvet går till den döda makens barn eller syskon.
Separat insamlat energiavfall ska packas i plastkasse eller papperspåsar.
Enligt Finlands lag ska alla människor behandlas likvärdigt.
Apotekfinska _ svenska
Österbottens TE-byråfinska _ svenska
Om du är studerande kan du söka en hyresbostad som är avsedd särskild för studerande.
I invånarhusen kan områdets invånare vistas och samlas samt få anvisningar och råd.
Finlands advokatförbundfinska _ svenska _ engelska
Volontärarbetefinska _ svenska _ engelska
Utkomststödet är avsett som en tillfällig hjälp.
En del universitetsstudier leder direkt till ett yrke.
Du kan också förbättra dina språkkunskaper.
Det är bäst att börja med en rutt som märkts ut.
Därför varierar även bidragens belopp och grunder.
Män och kvinnor badar bastu olika tider.
Vanda område har varit bebott länge.
Föräldrarna bestämmer barnets religion.
Telefon: 0800 414 004
Om du vistas i Finland tillfälligt, kan du få en finsk personbeteckning om det behövs till exempel på grund av ditt arbete.
Vanligen närvarar köparen och säljaren av bostaden samt bostadsförmedlaren, om en förmedlare har använts.
Flera olika Vi läser tillsammans-nätverk är verksamma på olika håll i Vanda.
Finländarna värdesätter också sin integritet och privatsfär.
Tolken är med på möten mellan dig och myndigheten.
Ingen får missgynnas på grund av dessa omständigheter.
Nupoli - hjälp för ungafinska _ svenska
Mer information om skilsmässa och upplösande av ett registrerat parförhållande hittar du på InfoFinlands sidor Skilsmässa.
Om du under en lång tid tar hand om ett sjukt eller handikappat barn under 16 år kan du söka specialvårdpenning (erityishoitoraha) från FPA.
Om du arbetar i Finland, kan du ha rätt till den offentliga hälso- och sjukvården även om du inte har en hemkommun i Finland.
Vård av barnet
Läs mer på Vanda kyrkliga samfällighets webbplats.
Med intyget kan du bevisa att du omfattas av den sociala tryggheten i Finland även om du arbetar utomlands.
Ungdomsgårdarna är öppna för alla ungdomar i åldrarna 9–17.
De 1–18 vardagar av faderskapsledigheten som du kan ta ut samtidigt med barnets mor kan delas upp i högst fyra perioder.
För unga under 30 år
Verksamhetsställen för handikappservicefinska _ engelska
Grundläggande utbildning.
Om du inte betalar en räkning eller en skuld, kan du få en betalningsanmärkning (maksuhäiriömerkintä) i kreditupplysningsregistret.
Befolkningen i Finland
020 634 0200 (på finska och på engelska)
Skyldigheter
Telefon: 0295 025 500
lör 9–15
Läs mer: Fritid.
På vissa orter finns det daghem, som fungerar på andra språk än finska eller svenska.
Hälsovård för högskolestuderandefinska _ svenska _ engelska
Öppet
Läs mer: Förlossning.
I Finland föder de flesta kvinnorna vaginalt.
Hushåll
Om du har antagits, meddela så fort som möjligt till läroanstalten att du tar emot studieplatsen.
Du kan också ta ut alla 54 faderskapspenningdagar separat, till exempel efter föräldraledigheten.
_ bulgariska
Du måste själv trygga din försörjning i Finland.
Alla finländska högskolor har ett eget stipendiesystem för de studerande som kommer från länder utanför EU/EES-området och som har godkänts för att avlägga en kandidat- eller magisterexamen på engelska.
Info om folkhögskolorfinska _ svenska
När hjälpbehovet är brådskande
Man får inte kräva sådana egenskaper av arbetssökanden som inte är nödvändiga i utförandet av arbetet.
Information om att ansöka studiestödfinska _ svenska _ engelska
När barnet har fötts
Om du har frågor om eller problem med din anställning, kan du kontakta anställningsrådgivningen för invandrare.
Om du är under 29 år gammal, bor i Vanda och inte har ett jobb eller en studieplats, kan du få råd och handledning i Kipinä.
Du kan även fråga om råd hos FPA.
Många människor flyttade från landsbygden till städerna och allt fler kvinnor började arbeta utanför hemmet.
Valmansföreningen ska ha minst 100 medlemmar.
Läs mer: Hyresbostad.
Konsumentskyddslagen (Kuluttajansuojalaki) tryggar konsumentens rättigheter i Finland.
Information om Hörselförbundetfinska
information om den sociala tryggheten och sociala förmåner
Klubbar
Vanligtvis får du en tidsfrist inom vilken du måste lämna Finland.
Befrielse från överlåtelseskatt på första bostadfinska _ svenska _ engelska
Att anmäla sig som arbetslös arbetssökandefinska _ svenska
Du kan delta i kurser under dagtid, på kvällar eller på veckoslut.
Du behöver en personbeteckning till för din arbetsgivare eller läroanstalt.
Därefter betalar du varje månad en bestämd summa det vill säga bruksvederlag (käyttövastike).
Var hittar jag jobb?
Kulturkonflikter hemma
En anställd vid TE-byrån tar kontakt med dig om det behövs ytterligare uppgifter.
Tidningar i Finlandfinska
Tänk på att privata hälso- och sjukvårdstjänster är avgiftsbelagda.
Du kan få behovsprövad rehabilitering om ditt mål är att fortsätta arbeta, återgå till arbetet eller börja arbeta.
Hjälptelefonen betjänar på många olika språk.
Staden och landskommunen slogs samman till nya Rovaniemi stad år 2006.
När finländare samtalar, kan det ibland uppstå tysta stunder.
Du får då din skattedeklaration till rätt adress.
Närmare beskrivningar av de olika färdighetsnivåerna finns på Utbildningsstyrelsens webbplats.
uppdrag inom vetenskap, kultur och konst
Av dem hör emellertid endast en del till de islamska samfunden.
Guide för arbets- och näringsbyråns invandrarkunder(pdf, 5,1 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ arabiska _ kurdiska _ thai _ vietnamesiska
Lär dig finska eller svenska
Information om fristående examenfinska _ svenska _ engelska
Du får kontakt med diskrimineringsombudsmannens byrå:
Skatteprocenten (Veroprosentti) beräknas i Finland för var och en separat.
Om en graviditet inte börjar inom ett år efter att man slutat använda preventivmedel kan saken undersökas.
Nämnden kan även stöda en förlikning mellan parterna.
Rådgivning tillhandahålls till exempel av:
När du flyttar till Finland måste du ansöka om uppehållstillstånd hos Migrationsverket eller registrera din uppehållsrätt.
Fastighetsförmedlingsbyråer och privatpersoner hyr ut bostäder även för korta perioder.
Vasa ortodoxa församlingfinska _ engelska _ ryska
Jobbsökning
I Helsingfors ordnas förskoleundervisning (esiopetus) i många daghem och skolor.
I förväg meddela till bostadsaktiebolagets disponent eller styrelse om du ska göra en sådan ändring i din bostad som kan påverka husets bärande konstruktioner, vattenledningar, fuktisolering, elledningar eller ventilationssystem.
Läs mer: Handikappade personer.
Läs mer på InfoFinlands sida Officiellt intyg över språkkunskaper.
Problem med uppehållstillståndet
Kurser i svenskafinska _ svenska _ engelska
Yrkesinriktad arbetskraftsutbildning är kostnadsfri.
Ett sätt att fira en helgdag är att hissa flaggan.
Om du ansöker om en plats i ett privat daghem, kontakta direkt det daghem som är föremål för platsansökan.
Barnet kan få uppehållstillstånd på grund av familjeband om hans/hennes förälder är finsk medborgare eller gift med en finsk medborgare och bor i Finland.
Information om att ansöka om arbetslöshetsersättning hittar du på InfoFinlands sida Arbetslöshetsförsäkring.
I Finland finns även privata mödrarådgivningar.
Du hittar mer information till exempel på Kehitysvammaliittos och Kehitysvammaisten Tukiliittos webbplatser.
Förskoleundervisningen börjar i augusti och ansökningstiden är i januari.
Avainboendefinska
Om ett barn blir sjukt under skoldagen vårdas han eller hon i skolan.
Hemvårdsstöd kan i vissa fall även betalas till familjemedlemmar som vistas i ett annat EU- eller EES-land.
Om makarna inte har upprättat ett äktenskapsförord, räknas båda parternas egendom med i bodelningen och egendomen delas jämnt mellan makarna.
Ohjaamo är en rådgivningstjänst som är avsedd för unga vuxna.
Vårdgarantifinska _ svenska
Om du behöver akut hjälp av tandläkaren på kvällen eller veckoslutet, ring jouren på tfn 09 471 71110.
Då kan sakerna som ligger på spisen fatta eld.
Barn kan ha fritt inträde till vissa museer.
Din situation avgör hur du kan finansiera dina studier i Finland.
Skyldighet att följa Finlands lagar även annanstans än i Finland.
Fråga mer om detta vid beskickningen för ditt eget land.
Hattulavägen 2
Den är en hälsosam och nästan gratis motionsform.
Rovaniemi karttjänstfinska _ svenska _ engelska
De kan få ett permanent uppehållstillstånd när äktenskapet har varat fem år.
I examen ingår olika uppgifter där följande färdigheter krävs:
Skicka din ansökan till adressen:
Om dina studier i Finland till exempel varar mindre än två år, ska försäkringen täcka sjukvårdskostnader upp till minst 120 000 euro.
Rättshjälpsbyrån i Rovaniemi
För varje studerande upprättas en personlig utvecklingsplan för kunnandet (PUK).
Biblioteket finns även på nätet.
Kom ihåg att skaffa eventuell flytthjälp i tid.
Grankulla hälsostation
I Finland råder religionsfrihet (uskonnonvapaus).
Även barnet måste vara närvarande när tillståndsansökan lämnas in.
Tillstånd och anmälan som är anknutna till idkandet av en näringfinska _ svenska _ engelska
Efter en preliminär undersökning får du en remiss till fortsatta undersökningar om det behövs.
Krismottagningen betjänar på finska, svenska och engelska samt på andra språk med hjälp av tolk.
Förberedande utbildning inför yrkesutbildning
Läs mer: Flytta till Finland.
Du får därför inget studiestöd (opintotuki) och inga studentrabatter när du studerar vid öppna högskolan.
I Finland är beskattningen progressiv.
Påsken är en kristen fest.
Finlands Röda Kors De ungas skyddshus (Suomen Punaisen Ristin Nuorten turvatalo) ger stöd och hjälp i krissituationer för 12–19-åringar.
Registerbeskrivning för InfoFinland finns på Helsingfors stads webbplats.
Skuldlinjen
Då du får en bostad ska du göra ett skriftligt bostadsrättsavtal (asumisoikeussopimus) med husets ägare.
Ofta använder man bedömningsskalan enligt den gemensamma europeiska referensramen (GER).
på svenska: 0295 020 711
Tjänsten är kostnadsfri för kunderna, dvs. du betalar endast din egen samtalskostnad.
Helsingfors stad har ett finskspråkigt arbetarinstitut och ett svenskspråkigt arbetarinstitut.
När du håller på att flytta till Finland, får du ytterligare information i avsnittet Flytta till Finland.
InfoFinlands chefredaktör och ansvariga redaktör är Eija Kyllönen-Saarnio.
Flerspråkiga biblioteketfinska _ svenska _ engelska _ ryska
Juristtjänsterna är avgiftsbelagda men om du har låg eller medelhög inkomst, kan du få gratis eller delvis ersättningsgill juridisk hjälp vid statens rättshjälpsbyrå (oikeusaputoimisto).
I hälsovården av 1–6-åriga barn får man hjälp av rådgivningsbyråns (neuvola) hälsovårdare och läkare.
Den viktigaste delen i affärsverksamhetsplanen är verksamhetsplanen för ditt eget företag.
I Sandudd finns dessutom Helsingfors ortodoxa begravningsplats, Helsingfors judiska begravningsplats och Helsingfors muslimska begravningsplats för tatarer.
Finnkino linkkiFinnkino:
Läs mer på InfoFinlands sida Boende för studerande.
I Helsingfors finns även några sådana gymnasieskolor där undervisningsspråket är något annat än finska eller svenska.
Information om den förberedande undervisningenfinska _ engelska
en hörselskada eller
linkkiRäddningsbranschens Centralorganisation i Finland:
Kartorfinska _ svenska _ engelska
Du har svenskspråkiga familjemedlemmar eller släktingar.
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Om du inte kan finska eller svenska kan du anlita en tolk när du sköter ärenden med myndigheter.
I annat fall betalar du en källskatt (lähdevero) på 35 % på lönen och du behöver ett källskattekort.
Självständighetsdagen
Vederlagen används till att sköta bostadsaktiebolaget, till exempel underhålla byggnaderna och gårdsområdet.
Du har även möjlighet att överklaga ett negativt beslut till förvaltningsdomstolen.
Du kan besöka vilket apotek som helst.
Olika företagsformer i Finland är firma, öppet bolag, kommanditbolag, aktiebolag och andelslag.
I den skrivs det in vilka studier du avlägger och hur.
Stadens befolkning växte snabbt och och på de inkorporerade områdena byggdes många nya förorter på 1950−1980-talen.
Finland är ett tvåspråkigt land
Stadsmuseetfinska _ svenska _ engelska
Till skillnad från äktenskap
uppfyller villkoren för inkomstrelaterad dagpenning, grunddagpenning eller arbetsmarknadsstöd.
Ett viktigt mål är att eleverna lär sig att tänka självständigt och tar eget ansvar för sitt lärande.
Tjänsten finns på finska, svenska, engelska, ryska, estniska, franska, somaliska, spanska, turkiska, kinesiska, persiska och arabiska. De olika språkversionerna är identiska.
Följande rättigheter och skyldigheter gäller även utlänningar bosatta i Finland.
Ni fattar gemensamt beslutet om på vilket sätt graviditeten avbryts.
Kommunens invånare har enligt kommunallagen rätt att lämna in motioner till kommunen i ärenden som gäller dess verksamhet.
Om du har kommit till Finland som kvotflykting har du hemkommun i Finland och rätt att utnyttja de offentliga hälsovårdstjänsterna.
Undervisning i finska för vuxna
Dessa tjänster hjälper människorna att klara sig bättre hemma.
Kontaktuppgifter till rådgivningsbyråerna
Dessa studier är vanligtvis avgiftsbelagda.
När du åker till sjukhuset ska du ta med dig tillräckligt varma kläder för barnet för hemresan.
Information om familjepensionfinska _ svenska _ engelska
Om din ledighet varar i 12 vardagar eller mindre, ska du meddela om ledigheten till din arbetsgivare en månad på förhand.
När du söker till en yrkesinriktad vuxenutbildning, ska du ha en tillräckligt lång arbetserfarenhet.
Du kan få arbetsmarknadsstöd om du
På en privat hälsostation måste kunden själv betala samtliga kostnader.
Om ett barn är i livsfara eller har hamnat i en olycka ska du ringa nödnumret (hätänumero) 112.
Om hyresavtalet kräver att du har en hemförsäkring, måste du teckna en sådan.
Vad innehåller ett CV?
tfn 040 152 3918.
Information om avfallshanteringfinska _ svenska _ engelska
Registrering av ett religiöst samfundfinska _ svenska _ engelska
Finland förklarade sig självständigt den 6 december 1917 och bolsjevikregeringen som tog makten i samband med oktoberrevolutionen i Ryssland erkände självständigheten den 31 december 1917.
Läs mer: Våld.
I Esbo finns motionsslingor och friluftsleder på olika håll i staden.
Om ärendet inte kan lösas på arbetsplatsen, ska du kontakta arbetarskyddsdistriktet (työsuojelupiiri) i ditt område eller ditt fackförbund.
Du hittar information om TE-byråns tjänster på InfoFinlands sida Om du blir arbetslös.
Om du är studerande kan du få en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS.
Arbete utan uppehållstillståndfinska _ svenska _ engelska
De ungas skyddshusfinska _ svenska _ engelska
Hur ansöker jag till yrkesinriktad arbetskraftsutbildning?
Anställningen ska vara minst fyra månader lång och din arbetstid och lön ska vara tillräcklig.
Också barn under 18 har rätt att fatta beslut i vissa ärenden.
I Finland ordnas stödboende (tukiasuminen) och serviceboende (palveluasuminen) för dem som behöver stöd för att kunna bo självständigt.
skriftliga färdigheter
Dessa uppgifter är till exempel namn, födelsedatum, nationalitet, kön och adress.
Du kan göra anmälan med ditt eget namn eller anonymt.
Intyget är giltigt i fyra månader.
linkkiExpatFinland.fi:
Mer information får du på Tullrådgivningen +358 (0)295 5201 eller på tullens webbplats.
Behovet av närståendevård bedöms inom seniorrådgivningen.
Om ditt företag är i förskottsuppbördsregistret kan du fakturera kunder utan förskottsinnehållning.
Som elevens egen religion undervisas bland annat islam, buddhism och ortodox religion, beroende på antalet elever.
Om du inte är säker på att isen håller, gå inte ut på isen.
Veckans bioprogram publiceras ofta också i lokaltidningen.
Det är också ett brott att föra en flicka till ett annat land, för att låta henne genomgå omskärelse där.
Läs mer: Sexualhälsa
Mer information om krävande medicinsk rehabilitering fås av FPA.
Om föräldrarna är gifta ska båda föräldrarna underteckna blanketten.
Familjen kan ändå söka rätt till småbarnspedagogik på heltid om barnet behöver särskilt stöd till exempel i att lära sig det finska språket eller på grund av att familjen befinner sig i en svår situation.
Socialarbetare 016-322 3126, 040-351 6925
När den unga har fullgjort sin läroplikt får han eller hon arbeta heltid mellan klockan 6.00 och 22.00.
FPA ordnar inte en annan tolk.
Idrottstjänsterfinska _ svenska _ engelska
Registrering av fordon på Internetfinska _ svenska _ engelska
Tolkcentralernas tjänster är främst avsedda för myndigheter som arbetar med invandrare.
Kurssökningen för kurser i finska och svenska, Finnishcourses.fi, är en del av InfoFinland.
I Finland får läkemedel inte säljas annanstans.
Fundera på vad arbetsgivaren bör veta om dina färdigheter och ditt kunnande.
Vailla vakinaista asuntoa ry. är en förening som hjälper bostadslösa.
Handikappbidrag för vuxnafinska _ svenska _ engelska
Avtalsparterna driver och utvecklar tjänsten tillsammans.
Fastlagen inleder förberedelserna för påsken.
Om du vill kan du även föda barnet på något annat sjukhus inom samkommunen Helsingfors och Nylands sjukvårdsdistrikt (HNS).
Då du köper ett egnahemshus köper du en fastighet.
Särskilda tjänster för utvecklingsstörda är bland annat
Du kan köpa tågbiljetter på VR:s webbplats, på järnvägsstationer och ombord på tågen.
Om du flyttar stadigvarande till Finland eller EES-området behöver du inte Patent- och registerstyrelsens tillstånd för att grunda företaget.
Du kan berätta vilka målsättningar du har med jobbsökningen eller vilken specialkompetens du besitter.
Vid RAMK finns det elva finskspråkiga och tre engelskspråkiga utbildningsprogram som leder till yrkeshögskoleexamen, fem utbildningsprogram som leder till högre
du är familjemedlem till en medborgare i ett EU-land, ett EES-land eller Schweiz
Den offentliga rättshjälpen finns även tillgänglig på engelska och vid behov kan man använda tolktjänster.
Vid Takuusäätiö kan du även ansöka om ett litet lån, om du behöver pengar för en utgift av engångskaraktär, såsom en hushållsmaskin, möbler, hyresdeposition, reparation av bilen eller glasögon.
Hyresbostad
linkkiBiblioteken.fi:
Du kan själv be om en inledande kartläggning.
Mottagande av studieplats
sambor
Du kan själv kontakta familjerådgivningen och komma överens om ett möte.
En del arbetsgivare ordnar undervisning i det finska språket för sina anställda.
Om du lämnar Finland under vistelsen och inte stannar i landet tre månader utan avbrott, behöver du inte ansöka om registrering av uppehållsrätten.
Terapi för unga kan också omfatta besök av föräldrar.
Du behöver ändå inte betala överlåtelseskatt om alla följande villkor uppfylls:
Om du vill grunda ett uppstartsföretag i Finland kan du ansöka om uppehållstillstånd för uppstartsföretagare som är avsett för tillväxtföretagare.
Familjen kan ansöka om utkomststöd om den har ekonomiska problem som den inte klarar av annars.
Länkar för frilansarefinska
MoniNetfinska _ engelska
Hos familjerådgivningen får barn, unga och familjer hjälp med problem som rör fostran av barn och barns utveckling.
Den unga har rätt att öppna ett eget bankkonto och förvalta de medel som han eller hon förtjänat med sitt eget arbete.
Om du har bokat tid, men inte kan komma, är det väldigt viktigt att du avbokar besöket i tid, vanligen senast dagen innan.
Efter det måste du förnya din ansökan om du fortfarande letar efter bostad.
linkkiRovala:
Vissa arbetsgivare ordnar finskundervisning för sina arbetstagare.
I vissa bostadsaktiebolag har man beslutat att fördela ansvaret på ett annat sätt.
Banker och Finnvera beviljar lån till företagare som startar ett företag.
Betala hyresgarantin senast på det datum som överenskommits i hyresavtalet.
Du behöver en skattenummer (veronumero), om du arbetar på en bygg- eller monteringsarbetsplats i Finland.
Finland är indelat i kommuner som har självstyre.
Tionde klasserna
Hälsostationerna har öppet mån–fre kl. 8.00–16.00.
I storstäderna kostar boendet mycket mer än på mindre orter.
Filmklipp om lekparksverksamhetfinska _ svenska _ engelska _ somaliska _ persiska _ arabiska
Du kan också anmäla dig till den inledande kartläggningen vid TE-byrån.
skattebyråerna,
I Finland tryggar lagen arbetstagarnas rätt att höra till ett fackförbund (ammattiliitto).
Ansökan om föräldradagpenningar
Hyresbostad.
På familjerådgivningscentralen får du hjälp om ni har problem i familjen eller i parförhållandet.
På långfredagen minns man Jesu död.
Efter gymnasiet kan man söka till universitet, yrkeshögskola eller gymnasiebaserad yrkesutbildning.
År 1972 fick köpingen stadsrättigheter.
De beslutar också huruvida dina utländska studier och din övriga kompetens kan godkännas som en del av den examen du avlägger i Finland.
linkkiKommunikationsverket:
Läs mer på InfoFinlands sida Fackförbund.
De övriga medlemskommunernas egna redaktioner upprätthåller sina egna kommunsidor.
Du kan köpa resekortet på Grankulla stadshus.
Grundläggande information om Finland
Kontaktuppgifterfinska _ engelska _ ryska _ franska _ arabiska _ rumänska _ bulgariska
Finska och svenska är Finlands nationalspråk.
Val i Finlandfinska _ svenska _ engelska
Språkkaféer:
Tips för jobbsökningenfinska _ svenska _ engelska
I Esbo beslutas ärenden av stadsfullmäktige.
Bifoga apotekets utredning över de köpta läkemedlen och kassakvittot.
Lapplands läroavtalscenter
Telefonnummer: 0295 025 500
Därför är det en tryggare boendeform än en ägarbostad.
En ny företagare får en rabatt på 22 procent på pensionspremierna under de fyra första åren.
Bifoga till din ansökan blanketten Boende och arbete utomlands.
Platsen för utförandet av arbetet
Om avtalet varit i kraft i kortare tid än ett år, är uppsägningstiden tre månader.
Besöksadress: Karlebygatan 27, 67100 Karleby
Mer information om den sociala tryggheten i Finland hittar du på FPA:s webbplats och på InfoFinlands sida Den sociala tryggheten i Finland.
Adress:
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
Grundläggande information om vigseln finns på magistratens webbplats.
När ett äktenskap slutar beslutar barnets föräldrar hur vårdnaden ska ordnas.
Hur länge man bor i stödbostad beror på kundens livssituation och behov.
Förskoleundervisningfinska _ svenska _ engelska
De integrationsrelaterade socialtjänsterna omfattar rådgivning och handledning.
Dessutom är en del av räntan på bostadslånet avdragsgill i beskattningen.
I detta fall avvisas du tillbaka till det land där du var innan du kom till Finland.
du inte är arbetslös, men du ska gå över till företagande på heltid till exempel från lönearbete, studier eller arbete i hemmet.
Kontaktuppgifter till De ungas skyddshus:
Länderna som tillhör Schengenområdet har enhetlig visering.
På yrkeshögskolan är undervisningen mer praktiknära än på universitetet.
Vuxenutbildningsinstitutet ligger i Dickursby, men kurser ordnas runtom i Vanda.
I lagstiftningen och kollektivavtalen fastställs till exempel minimilöner, arbetstider, semester, lön under sjukskrivning och uppsägningsvillkor.
I Finland kan kvinnor och män själva besluta vem de ska gifta sig med.
om hur du kan återhämta dig.
Blanketten får du antingen vid informationen på Grankulla stadshus, på socialbyrån eller på Grankulla stads webbplats.
Rådgivningarna för familjeplaneringfinska _ svenska.
tfn 010 8022 40
Vanligtvis går det inte att få tag på en tolk snabbare än så.
Info om sommaruniversitetfinska _ svenska
Kommunen kan även ge dig servicesedlar med vilka du kan köpa tjänsten av en serviceproducent som kommunen godkänt.
Spiralen passar bäst för kvinnor som har fött barn.
Syftet med projektet är att utveckla tjänsteprocesserna för invandrare, avsedda för den inledande tiden direkt efter inflyttningen.
AA-grupper finns på många orter och i de större städerna finns även grupper på engelska.
Läs mer om handikappbidrag för barn och specialvårdpenning på InfoFinlands sida Ett handikappat barn.
Via det kan du få en mentor som stöder dig när du söker arbete eller studieplats eller grundar ett företag.
En myndighet, till exempel en notaries publicus, måste verifiera överenskommelsen.
Till exempel mat och många typer av tjänster kostar i genomsnitt mer i Finland än i övriga Europa.
Du kan söka skilsmässa ensam eller tillsammans med din maka/make.
Oy
Om du är i Finland som turist och råkar ut för någon besvärlig situation, kontakta ditt hemlands beskickning.
du har varit fortlöpande bosatt i Finland under minst ett års tid.
Olika företagsformer i Finland är enskild näringsidkare (toiminimi); öppet bolag (avoin yhtiö); kommanditbolag (kommandiittiyhtiö); aktiebolag (osakeyhtiö) och andelslag (osuuskunta).
Ett arbetsavtal uppstår när arbetstagaren och arbetsgivaren kommer överens om utförandet av ett arbete och lönen som betalas för det samt övriga förmåner och villkor.
Det finländska sättet att kommunicera är rakt och okomplicerat.
Det är bra att ta reda på hur stora lönerna är i den egna branschen i Finland.
Jämlikhet inom hälsovården
du har fått humanitärt skydd, men ditt uppehållstillstånd löper ut eller har redan löpt ut.
I Finland utgörs en familj av
Läs mer: Bostadslöshet.
I Finland finns sex regionförvaltningsverk.
Det är viktigt att sätta upp tydliga gränser och regler för barn och unga.
Om du flyttar till en kommun där ditt bibliotekskort inte gäller, måste du skaffa dig ett nytt bibliotekskort vid biblioteket på din nya hemort.
någon är i livsfara (hengenvaara)
Om du behöver juristens hjälp med något som har med uppehållstillstånd eller ansökan om finskt medborgarskap att göra kan du kontakta Flyktingrådgivningen som har jurister specialiserade på tillståndsärenden.
Planera noga
Läs mer om myndiga medborgares rättigheter och skyldigheter på InfoFinlands sida Dina rättigheter och skyldigheter i Finland.
Anmälan till hemspråksundervisning görs varje år i mars.
inte är gifta eller under förmynderskap.
företagande som huvudsyssla
Finlands ställning under självständighetens tidiga år var skör.
Du kan också studera vid en yrkesläroanstalt och ett gymnasium samtidigt.
Om pojken är gammal nog för att säga sin åsikt ska han tillfrågas om han samtycker till operationen.
Du kan använda en tolk när du vill om du beställer tolken själv och betalar kostnaderna.
Lapplands läroavtalscenterfinska
Om ordföranden eller vice ordföranden har sin hemort utomlands kan föreningen ansöka om dispens hos patent- och registerstyrelsen.
Det finns många bussbolag i Finland.
du är intresserad av högskolestudier och
Ansökan till universitetfinska _ svenska _ engelska
Mer information finns på InfoFinlands sida Hemkommun i Finland .
Försäkrings- och finansrådgivningen
På De ungas skyddshus kan du få samtalshjälp och tillfällig logi.
I stadens skolor är undervisningsspråket finska eller svenska.
Kärnkraftverket levereras av RAOS Project Oy, ett bolag som ingår i den ryska Rosatom-koncernen.
De är finsk-ugriska språk.
Socialjouren (sosiaalipäivystys) hjälper kvällstid och under veckoslut om du är i akut behov av hjälp av en socialarbetare.
Grankulla är en av de fyra kommunerna i huvudstadsregionen.
För frågor gällande jouren ring tel. (06) 828 7450.
Om du köper en fastighet är skatten 4 procent av bostadens skuldfria pris.
Föreningen för familjer med en förälder (Yhden Vanhemman Perheiden Liitto) ger information och ordnar aktiviteter för familjer med en förälder.
FPA ordnar yrkesinriktad rehabilitering för unga personer och vuxna som inte arbetar.
Karleby familjerådgivning
Seniorrådgivningenfinska _ svenska
Brådskande tandvård/första hjälpen (nattjour):
Öppet varje dag kl. 17–10.
Information om CVfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
Det kan vara svårt att hitta en bostad med lämplig hyra.
Båda makarna måste vara på plats vid vigseltillfället.
Om du flyttar till Finland för att arbeta från EU-området eller ett EES-land eller Schweiz, omfattas du vanligtvis av den sociala tryggheten i Finland under din anställning, även när din anställning är kortvarig.
Du kan fylla i ansökan på Internet eller posta den till FPA.
Ansökan om Karleby stads hyresbostadfinska _ svenska _ engelska
Intyg över äktenskap eller registrerat parförhållande
linkkiOhjaamo:
Finlands folkmängd är cirka 5,5 miljoner människor.
Hyresgästens rättigheter och skyldigheter
Hem och familjsvenska _ engelska _ ryska _ estniska
Du kan också ansöka om oavlönad ledighet om din situation kräver att du är frånvarande en längre tid.
Information om Konstskolanfinska _ svenska
dickursbyvägen 44 F, vån.
I Esbo finns flera rådgivningsbyråer på olika håll i staden.
En jobbansökan är oftast en knapp sida.
Dina familjeförhållanden och andra kontinuerliga pensionsinkomster påverkar också folkpensionens belopp.
Om du vill träffa en kvinnlig läkare, ange detta när du bokar tiden.
Du kan påvisa dina språkkunskaper:
En ny företagare kan anmäla sig till Skatteförvaltningens förskottsuppbördsregister.
Den viktigaste lagen är grundlagen( perustuslaki).
Det lönar sig att jämföra kommunalt ägda och privata servicehus.
Frivilligarbete är oavlönat arbete, men arbetserfarenheten kan vara nyttig när du söker ett avlönat arbete.
I karttjänsten visas även var största delen av motionsplatserna finns.
Om du blir utsatt för ett brott, gör en brottsanmälan hos polisen.
Rautbergsgatan 3
En utredning över att ni har bott tillsammans i två år eller har gemensam vårdnad om ett barn, om du är i ett samboförhållande
Du hittar närmare information i Studieinfo.fi.
När du blir sjuk ska du först kontakta din egen hälsostation (terveysasema). Där kan du boka tid hos en allmänläkare eller en hälsovårdare.
Europeiska recept kan skrivas ut av yrkesutbildade personer inom hälso- och sjukvården som arbetar i ett EU- eller EES-land eller Schweiz och har förskrivningsrätt.
Alla bibliotek har en webbplats där du kan söka information om bibliotekets samlingar och förnya dina lån samt reservera material.
Ett tidsbestämt hyresavtal kan inte sägas upp mitt i avtalsperioden.
Man får syskonrabatt.
Under kvällar och veckoslut finns jourmottagningen för barn under 16 år vid Jorv sjukhus och på Barnkliniken i Helsingfors.
polisen,
Denna regel gäller till exempel utbytesstudenter som endast studerar en kort period i Finland (t.ex. fyra månader). Om du lämnar
Pensionssystemet i Finlandfinska _ svenska _ engelska
Under tiden då din ansökan behandlas kan du få rådgivning och rättshjälp vid den offentliga rättshjälpsbyrån.
Skattekort och skattenummer
Social- och hälsostationen i Kilo
FPA kan betala ut understöd för psykoterapin, men du måste själv hitta en lämplig terapeut.
En väsentlig del av studierna är inlärning på arbetsplatsen.
De övriga är hembygdsmuseer som vanligen bara har öppet sommartid.
Nätstöd för ungdomar, Nuortennettifinska
Fpa ersätter arbetsgivaren och företagaren en del av kostnaderna för företagshälsovården, om dessa är nödvändiga och rimliga.
Minst 20 myndiga personer kan grunda ett religiöst samfund.
I en krissituation kan du ringa nödcentralen på numret 112.
Läs mer: Stöd för vård av barn i hemmet
linkkiFlyktingrådgivningen rf:
På vintern fryser de flesta vattendrag till i Finland.
Sökning av ägarbostäderfinska _ engelska
moderskapsledighet
I den finländska arbetskulturen tilltalar man varandra på ett mycket informellt sätt.
Om du besöker jouren kvällstid eller under helger ska du först ringa jourens telefonrådgivning (06) 826 4500.
När du gifter dig kan du
Med hjälp av menyn Städer får du fram information om den kommun som du är intresserad av.
Hilma för handikappade invandrare som erbjuder servicevägledning och rådgivning för handikappade invandrare och långtidssjuka.
Fackförbundet och arbetslöshetskassan är dock två separata system.
när den ena makan eller båda makarna tillsammans kräver att de ska dömas till skilsmässa.
Den största av dem är Helsingfors-Vanda flygplats.
De erbjuder även mycket nyttig information och tjänster till hörselskadade.
Du kan vara offer för människohandel, om
Telefon: (06) 8287 580
Krävande medicinsk rehabiliteringfinska _ svenska _ engelska
Det kan till exempel vara vardagliga tips om arbete, studier, tillståndsärenden, boende eller språkinlärning.
Karleby blev en viktig industristad främst tack vare läder- och metallindustrin.
Det finns även hemlika lägenhetshotell med lägenheter som till exempel kan ha ett eget kök.
Om barnets förälder har uppehållstillstånd på grund av internetionellt skydd, men inte flyktingstatus, krävs att föräldern har en tillräcklig inkomst för att barnet ska kunna få uppehållstillstånd.
Barnkapningar (lapsikaappaus)
Fråga mer vid din egen hälsostation under dess öppettider eller leta upp informationen på din hemkommuns webbplats.
Läs mer: Behöver du en jurist?
Alexandersgatan 9, 4:e våningen (Köpcentret Kluuvi)
Äktenskap.
på en blankett som du får på posten eller hos magistraten.
Anställda inom företagshälsovården har sekretessplikt.
Vid mödrarådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Förbundet strävar efter att trygga sina medlemmars intressen i arbetslivet.
Du kan ansöka om folkpension om du inte har någon arbetspension eller om din arbetspension är väldigt liten. Folkpensionens belopp beror på hur länge du har bott eller arbetat i Finland.
Detta hjälper om det uppstår konflikter i arbetet.
Namnlagenfinska _ svenska
Förlåt.
Högskolor ordnar engelskspråkig undervisning i vissa utbildningsprogram.
Småbarnspedagogik är fostran, undervisning och omsorg som är pedagogiskt planerad och som har noga genomtänkta mål.
Övrigt kunnande – Språkkunskaper, IT-kunskaper, avlagda tillståndskort, till exempel hygienpass.
Handikappade personerlinkkiEsbo stad:
En del appar kostar pengar.
Parktanterfinska
som inte står under förmyndarskap
Vid problem i parförhållandet kan du söka hjälp till exempel vid familjerådgivningen eller hälsovårdscentralen i din hemkommun.
Om du inte har betalat en räkning senast på förfallodagen får du en betalningspåminnelse.
Du kan få tillståndet om:
Mor- eller farföräldrarna bildar en egen familj.
Du kan också få blanketten hemskickad per post.
Rådgivningsbyråerfinska _ svenska _ engelska
Arbetsavtalet är bindande för båda parterna.
Arbetsgivaren och arbetstagaren kan ändå i arbetsavtalet komma överens om villkor som är bättre än villkoren i kollektivavtalet.
Barnets underhållsbehov delas mellan föräldrarna enligt deras underhållsförmåga.
MIELI rf:s kristelefon erbjuder omedelbar samtalshjälp för människor i kris och deras närstående.
Moderskapsunderstödet är antingen en moderskapsförpackning (äitiyspakkaus) eller ett fast skattefritt belopp, du väljer vilket alternativ du vill ha.
Tolken ska vara vuxen.
Enligt Finlands lag får en människa inte diskrimineras på grund av sin sexuella läggning.
förföljelse och diskriminering
födelseattester för dina barn
Oyfinska
Du har rätt
Arbetslöshetsförmånerna är den inkomstrelaterade dagpenningen, grunddagpenningen och arbetsmarknadsstödet.
Du kan också komma överens med personalen om att din språkkunniga make eller vän tolkar under förlossningen.
självständighetsdagen 6.12
Hur skaffar jag en hyresbostad?
Du kan också fråga direkt vid läroanstalterna.
statlig tjänsteman
B2 – ASE 4
tfn 0400 187 250
Du ska aldrig placera något ovanför bastuugnen, använda bastun som förråd eller torka tvätt i bastun, eftersom detta kan orsaka en brand.
Information om hälsovården för skolbarnfinska _ svenska _ engelska
Medborgarinstitut
Hjälp med att söka jobb
Om du inte har hemvist inom EES och är medborgare i något annat land än ett medlemsland i den Europeiska unionen, ett EES-land eller Schweiz, behöver du ett uppehållstillstånd för att driva ett företag i Finland.
Pensionsförsäkringar fås antingen genom försäkringsbolag eller pensionskassor (eläkekassa).
Läs mer om föräldrarnas skyldigheter gentemot sina barn på InfoFinlands sida Fostran av barn i Finland.
Socialbyrån kan ha olika namn i olika kommuner.
Folkhögskolan kan drivas av en organisation eller också kan de vara självständiga institut.
Läs mer på InfoFinlands sida Hyresavtal.
Vandainfo ger dig information om såväl Vandas stads som statens tjänster.
Där kan man tala om problem och få hjälp och stöd.
Maria Akatemia hjälper kvinnor som har utövat våld eller fruktar att de kommer att utöva våld mot en familjemedlem.
Offentliga hälsovårdstjänster tillhandahålls vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
När socialväsendet bekräftar avtalet är det lika officiellt som ett domstolsbeslut.
Du kan även kontakta Kriscentret Monika via chatten.
På mödrarådgivningen och på vissa förlossningssjukhus ordnas familjeträning som ska hjälpa modern och familjen att förbereda sig för den kommande förlossningen och att ta hand om babyn.
Då måste du vänta på behandlingen av besvären utomlands.
God morgon!
Om barnet har fyllt tolv år måste man få barnets skriftliga tillstånd för att byta barnets efternamn.
Tfn 0800 05058
En välhållen bil kostar flera tusen euro.
Videoklippet ska vara i enlighet med Finlands lag och följa god sed.
Tjänsten är avsedd för män som flyttat till Finland, oberoende av bostadsort.
I svenskan böjs verben i olika tempus.
Till exempel på fester serveras det nästan alltid kaffe.
Invånarna i Vanda kan påverka beslutsfattandet och beredning av ärenden på många olika sätt.
Elevens närskola bestäms enligt gränserna för dessa områden. Närskolan är i regel den skola som ligger närmast elevens hem.
arbetarskydd
Riksomfattande föreningar för invandrare
Endast kvotflyktingar kan få ersättning för familjemedlemmarnas resekostnader.
Fråga om studier i svenska hos utbildningsväsendet i din hemkommun, studievägledarna vid läroanstalter eller rådgivningstjänsterna för invandrare.
Barnrådgivningarfinska _ svenska
Vem är berättigad till utkomstskydd för arbetslösa?
Esbo och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
Skicka din ansökan till Fpa:s byrå eller skicka in den på internet.
linkkiCentria yrkeshögskola:
linkkiFöretagsEsbo:
Om familjen får tvillingar är föräldrapenningperioden 60 vardagar längre.
Observera att hindersprövningen kan ta flera veckor om den kräver intyg från andra länder.
linkkiUtbildningsstyrelsen :
graviditeten varat i cirka fem månader
Du ansöker om studieplats direkt vid läroanstalten.
motion
Religionsfrihetfinska _ svenska _ engelska
Seniorrådgivningen bedömer behovet av anhörigvård för en äldre person.
I Finland finns det olika tjänster som främjar din integration, hjälper dig att hitta sysselsättning och lära dig språket.
I allmänhet ska dessa avgifter betalas direkt till husbolaget.
På fastlagen åker man i Finland backe och äter fastlagsbullar som har bland annat grädde som fyllning.
Beloppet som krävs ska finnas på ditt bankkonto eller också ska du ha ett intyg över ett stipendium som beviljats av en officiell instans.
Ny företagsverksamhet ska anmälas till handelsregistret som upprätthålls av Patent- och registerstyrelsen (Patentti- ja rekisterihallitus).
Vissa brottmål kan behandlas skriftligt i domstolen, och då behöver man inte delta i rättegången.
Många finländare uppskattar anspråkslöshet.
Du kan ringa Omatila-tjänsten dygnet runt. Du behöver inte uppge ditt namn när du ringer.
Kandidater kan nomineras av
Årliga helger
Bildningscentralen
Mathjälp och inkvartering
Om du vill ha rådgivning på engelska, ska du skicka in din fråga via Företagsfinlands engelskspråkiga webbplats.
Vid behov skriver läkaren en remiss till närmare undersökningar.
Så länge handläggningen av din första ansökan om uppehållstillstånd pågår har du inte rätt att arbeta.
Om familjens pengar inte räcker till att betala hyran för bostaden eller kostnaderna för en ägarbostad kan familjen ansöka om allmänt bostadsbidrag vid Fpa.
Du kan krävas på vårdkostnaderna i efterhand.
Det beror på din arbets- eller studieplats vilken examensnivå du måste avlägga.
Mer information om giftermål i Finland hittar du på InfoFinlands sida Ingående av äktenskap i Finland, komihåglista.
Observera att tävlingsdeltagaren ansvarar för att verket eller en del av verket, till exempel musik eller bilder, som skickas till tävlingen inte gör intrång på en tredje parts upphovsrätt, varumärkesrätt eller immateriella rättighet.
ett barn som förts utomlands inte har lämnats tillbaka till Finland vid avtalad tidpunkt.
JA: hemmets stora och små batterier, mobiltelefonens batteri
Jämlikhet
Tillståndet är alltså inte kopplat till din nationalitet utan till var du har din hemvist.
Om du har frågor om tjänsterna vid Grankulla stad kan du kontakta stadens rådgivningstjänst via e-post på adressen neuvontapalvelu(at)kauniainen.fi.
Enskild näringsidkare (toiminimi)
I Grankulla finns också ett engelskspråkigt daghem.
du är 18–39 år gammal
Utbildningsavtalet är inlärning i arbetet.
Du kan ansöka om faderskapspenning även om du är till exempel företagare, arbetslös eller studerande.
Rådgivning på engelska om beskattningen i Finland: 029 497 050
Domus Arctica-stiftelsens webbplatsfinska _ engelska
Hälsovård för invandrare och asylsökande
Biblioteket ligger i Böle i Helsingfors.
När du får uppehållstillstånd eller registrerar din uppehållsrätt, får du samtidigt skriftlig information om
I förskolan lär sig barnen bland annat matematik, miljö- och naturkunskap samt konst och kultur.
Lapplands yrkesinstitut erbjuder förberedande utbildning för invandrare som vill söka till yrkesutbildning.
I Esbo finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
Betala hyresdepositionen först när du har ett skriftligt hyresavtal.
Flerfaldigt medborgarskap kan vara en fördel, men också en nackdel.
Sändaren ska inhämta skriftliga tillstånd för framställning av videoklippet och för tillverkning av kopior av samtliga personer som medverkat i framställningen av videoklippet.
tel. 044 730 7640
1906 Allmän och lika rösträtt, även för kvinnor
I en sådan situation är det viktigt att man skaffar sig hjälp.
Sök till gymnasiet i den gemensamma ansökan till andra stadiet.
Magistraten i Helsingfors
På internet finns många bostadsförsäljningsannonser. Bostäderna i Esbo är tämligen dyra.
En företagare och andra som arbetar åt sig själv kan ordna företagshälsovård för sig själv om de så önskar.
Hjälp vid drogproblemfinska _ svenska _ engelska
Skriv en ny ansökan och uppdatera ditt CV varje gång när du ansöker om ett nytt jobb.
I Karleby finns flera olika religiösa samfund.
När du vårdar en närstående i hemmet
Vi tar gärna emot respons på och utvecklingsidéer med koppling till InfoFinlands verksamhet, översättningarna och samarbetsmöjligheter.
Metallen i batterierna årervinns och de farliga ämnena hanteras på ett säkert sätt.
Ett barn med en svår sjukdom eller ett handikapp kan även få FPA:s handikappbidrag för barn under 16 år (alle 16-vuotiaan vammaistuki).
Miehen Linja (Miehen Linja) är en tjänst som hjälper män, som har utsatt sina familjemedlemmar för våld. Tjänsten är avsedd för invandrarmän.
Du ska bifoga ett studieregisterutdrag till din ansökan om fortsatt uppehållstillstånd.
Under sommaren är det möjligt att repetera gymnasiestudier vid sommaruniversitetet.
De separata ansökningarna kan ordnas under olika tidsperioder och ansökningsförfarandena kan avvika från varandra.
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i servicehus (palvelutalo) eller på en vårdinrättning (laitos).
Friluftskartafinska
Bostadsrättsbostäder är inte förknippade med ekonomiska risker.
Att ansöka om skilsmässafinska _ svenska _ engelska
Unescos världsarv
Du kan ansöka om FPA:s åldringspension och garantipension även per telefon.
När du vill grunda ett företag ska du noga fundera på om du har en bra affärsidé.
linkkiPensionsskyddscentralen:
Barnskyddet stöder familjen även då ett barn eller en ung till exempel använder mycket rusmedel eller begår brott.
Du besöker arbetsplatser och deltar i verkstäder.
Invånarlokalen i Kivenkolo
Ett skriftligt avtal om de centrala villkoren i arbetet
Om du fått uppehållstillstånd och din hemkommun finns i Finland kan du använda tjänsterna inom den offentliga hälsovården på samma sätt som de övriga invånarna i kommunen.
Du kan även föra barnet till en privat läkarstation.
arbetsersättning
En företagare är arbetslös när han eller hon har lagt ned sin företagsverksamhet eller sålt sin andel av företaget.
Om ditt barn är i en psykiskt påfrestande situation kan du kontakta familjerådgivningen (perheneuvola) i din hemkommun.
Om du vill kan du ansluta dig till fackförbundet i din egen bransch.
Du kan anmäla dig som kund vid TE-byrån antingen vid den lokala TE-byrån eller på TE-byråns webbplats.
Skriv ansökan och CV på samma språk som används i annonsen.
Familjerådgivningen
Om en av föräldrarna vill sköta barnet hemma efter föräldrapenningperioden, kan han eller hon få hemvårdsstöd.
Skolan börjar i augusti och slutar i slutet av maj eller i början av juni.
Till exempel A-tulkkaus förmedlar i Helsingforsregionen kontakttolkar för tillfällen där du uträttar ärenden hos myndigheter.
Du kan även skriva ut anmälningsblanketten på nätet och lämna in den till polisstationen.
Familjerådgivningfinska _ svenska
Karleby är en kulturstad med mycket att se och uppleva.
linkkiVanda ekonomi- och skuldrådgivning:
Till exempel Noux nationalpark ligger delvis på Esbos område.
Om du har betalat för mycket i skatt, får du skatteåterbäring (veronpalautus).
Om familjen bor nära gränsen till Helsingfors eller Esbo, kan du också söka dagvårdsplats i grannkommunen.
Alternativen är fler på våren.
medborgarskap,
Motionsmöjligheterfinska _ svenska
Professionellt erkännande och rätt till yrkesutövning
När ska jag söka hjälp?
Du kan till exempel beställa ett nytt skattekort om du ha nätbankskoder eller ett mobilcertifikat.
Också kommunerna ordnar aktiviteter för barn och unga.
Du hittar kontaktuppgifterna till rådgivningen på Brottsofferjourens webbplats.
Ledamöterna i kommunfullmäktige, eller bara kommunfullmäktige, utses i kommunalval.
För detta fastställs en bassjälvrisk.
I affärsverksamhetsplanen funderar du på styrkorna och svagheterna i ditt kunnande och egenskaperna hos den produkt, vara eller tjänst som du erbjuder.
1640 I Åbo grundas
Jourmottagning för barnfinska _ svenska _ engelska
tfn 040 4873 010
NewCo Yritys Helsinki erbjuder individuell rådgivning om grundande av företag samt ordnar informationsmöten och företagarutbildning på flera olika språk.
Stöd med jobbsökningen för under 30-åringar vid Navigatorn
Traditionella minoriteter i Finland är till exempel finlandssvenskarna, samerna, romerna, judarna och tatarerna.
Om du flyttar till Finland för att bo här stadigvarande ska du också registrera dig som invånare i magistraten (maistraatti).
Mer information om språkcaféerna får du från biblioteken.
Också de personer som inte har rätt till den offentliga hälsovården i Finland kan besöka privata hälsostationer.
Utlåtandet ger dig dock inte kvalifikationer att utöva ett reglerat yrke i Finland.
Under andra världskriget kämpade Finland två krig mot Sovjetunionen: först vinterkriget åren 1939–1940 och därefter fortsättningskriget åren 1941–1944.
Den förberedande undervisningen förbereder barnet inför grundskolan.
Godtagbara orsaker för uppsägning definieras i arbetsavtalslagen.
Hjälp vid sexuellt våld
På andelslagets stämma har varje medlem en röst. Medlemmarna ansvarar för andelslagets förpliktelser (till exempel skulder) endast med det belopp som de investerat i andelslaget.
Till exempel föreningen för handikappidrott och -motion i Finland, VAU ry, ordnar olika idrotts- och motionsevenemang.
Den varmaste månaden är juli, då stiger temperaturen dagtid ofta över 20 grader.
Vem som helst kan studera vid de öppna högskolorna.
Barnets flerfaldiga medborgarskap
Rovaniemis färger bär ett budskap för övriga Finland och Europa om de anpassningsbara nordliga breddgraderna, den arktiska kulturen och människorna.
Polisen kan förlänga uppehållstiden för ditt visum eller visumets utgångstid om du av motiverade skäl inte kan lämna Finland när ditt visum utgår.
Företagsrådgivare
Du kan beviljas EU-uppehållstillstånd (P-EU) för tredjelandsmedborgare om:
Om du är EU-medborgare kan du ansöka om personbeteckning samtidigt som du ansöker om registrering av uppehållsrätt.
I mataffären säljs endast milda alkoholdrycker.
Partnern kan delta i beslutsfattandet om kvinnan vill ta hänsyn till hans åsikt.
Karleby stad erbjuder gratis förskoleundervisning för alla 6 år fyllda barn.
Bosättningen utvecklades först vid vattendrag och det finländska territoriet har alltid använts för livlig handelstrafik.
Flyttjänsterfinska _ svenska _ engelska
På den här sidan finns mer information om den finländska arbetskulturen.
Om du har din hemkommun i Vanda, kan du utnyttja de offentliga hälsovårdstjänsterna.
Presidentvalet har vanligen två steg.
samhälleliga områden
Du måste också anmäla dig till rösträttsregistret i Finland.
Ansökan om dagvårdsplatsfinska
Om föräldern har fått flyktingstatus den 1.7.2016 eller senare, ska man ansöka om uppehållstillstånd för barnet inom tre månader från att föräldern fått flyktingstatus.
Låt alltid barnets intressen gå först när ni beslutar om boendet.
Ambulanser är endast avsedda för allvarliga och brådskande situationer.
Det lönar sig att ansöka om bostad på flera ställen.
Innan du ansöker om pension ska du begära ett arbetspensionsutdrag av din pensionsanstalt eller Pensionsskyddscentralen.
Flyktingrådgivningen r.f.
I Esbo finns tre biografer.
Unga som saknar studieplats eller arbete kan få hjälp av det uppsökande ungdomsarbetet.
Information om posttraumatiskt stressyndromfinska _ engelska _ ryska _ franska _ somaliska _ turkiska _ persiska _ arabiska _ kurdiska _ albanska _ vietnamesiska _ burmesiska _ bosniska _ serbiska _ swahili
Särdrag i undervisningen
Du kan fråga om den grundläggande utbildningen och om skolorna i Helsingfors vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning.
En bostadsvisning ordnas oftast för alla intresserade på samma gång.
Vanligen har man en kort kaffepaus på förmiddagen, en lunchpaus mitt på dagen och en kaffepaus till på eftermiddagen.
Först efter detta registreras ditt barn i befolkningsdatasystemet.
Om barnet har ett annat modersmål än finska eller svenska, får hen stöd i lärandet av finska eller svenska.
Broschyr Information om äktenskapslagenfinska _ svenska _ engelska _ ryska _ arabiska
I januari 1918 tog det röda gardet, som representerade arbetarna, makten i HelsingforsHels.
Mottagning för unga finns vid Nupoli.
Du kan också kontakta arbetsgivaren och begära mer information, om du undrar över något som inte framgår av jobbannonsen.
Information för närståendevårdare(pdf, MB)finska _ engelska _ ryska _ somaliska _ kinesiska _ persiska _ arabiska _ kurdiska
Stadigvarande boende kan påvisas till exempel genom följande omständigheter:
Du kan ringa en arbetsgivare direkt eller skicka en öppen ansökan via e-post.
Rehabilitering för barn
Den kan också göras på ett annat ställe, t.ex. vid en läroinrättning.
Om du beställer en ny specifikationsdel, tas det ut en avgift för den.
Bifoga även till ansökan om uppehållstillstånd din egen redovisning av situationen.
Mötesspråket är engelska.
Du kan ansöka om rehabilitering vid arbetspensionsanstalten om du har arbetat fem år eller längre.
Införsel av bil till Finland som flyttsak
Om du på förhand vet att du behöver bostaden enbart för en viss tid, är ett tidsbestämt hyresavtal ett bra alternativ.
Efter föräldraledigheten kan barnet börja i dagvård eller någondera av föräldrarna kan vårda barnet hemma.
Bastun är en viktig del av den finländska kulturen.
Ansök om tillståndet i ditt hemland eller i ett annat land där du vistas lagligt.
Om du är medborgare i något av de nordiska länderna, ett EU-land, ett EES-land eller i Schweiz och kommer till Finland för att arbeta eller driva ett företag, måste du registrera din uppehållsrätt.
p. 050-597 1122
Information om fisketillståndfinska _ svenska _ engelska
Många flyttade till Finland även för att studera, arbeta eller för att de hade sin familj här.
Organisationens verksamhet i Finland omfattar informering, utbildning och socialarbete.
De är även lämpliga för studier i det finska språket.
Du kan söka information om rutterna i Reseplaneraren (Reittiopas).
Information om hobbymöjligheter för ungdomarfinska
Pojken har rätt att vägra att gå med på operationen.
linkkiBio Grani:
Storkisbackens tandklinik
Vetenskaplig fortbildning vid universitet är examensinriktad fortbildning.
Om endera parten hör till den evangelisk-lutherska kyrkan eller ortodoxa kyrkan kan ni också begära hindersprövning i den egna församlingen.
Tänk också på vilka produktionsmedel eller hurudan arbetskraft du behöver.
Arbetsgivaren drar av arbetstagarens andel från lönen och betalar den och sin egen andel av försäkringspremierna till pensionsanstalten.
Du behöver dock tillstånd till detta av husets ägare.
De kan till exempel hjälpa dig om du har råkat ut för en olycka, blivit sjuk eller fallit offer för ett brott.
arbetslöshetsdagpenning
du är misstänkt för ett brott som är belagt med fängelsestraff
Använd inte material, såsom bakgrundsmusik eller bilder, som en tredje part har upphovsrätt till.
Äktenskap som ingåtts utomlands
Om du blir bostadslös på grund av en kris eller en olycka, ska du kontakta socialbyrån.
Om du har barn och går igenom en skilsmässa ska du ta kontakt med barnatillsyningsmannen.
De behöver inte ha föräldrarnas tillstånd.
Du kan komma till *Lapplands mödra- och skyddshem om någon i din familj är våldsam eller om du på grund av hot om våld inte vågar stanna hemma.
Läs mer: Handikappade personer.
linkkiHelsingforsregionens miljötjänster:
Många finländare är kristna men inte speciellt religiösa.
Att lämna asylansökan utan prövningfinska _ svenska _ engelska
Äldre människor
Ansökan till universitet
Där får du hjälp när du söker bostad eller tillfällig inkvartering.
Många firar också med mousserande vin.
En registrerad förening kan ansöka om finansiering och bidrag samt samarbeta med andra föreningar och myndigheter.
Oftast bor man i heminkvartering ett par dygn eller veckor.
När du går till magistraten ska du ta med dig
Anvisning för identifiering av bröstcancer(pdf, 440kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ thai _ rumänska _ samiska
På separat överenskommelse kan vigseln också förrättas någon annanstans, till exempel hemma eller i en festlokal.
Du kan även fråga om andra saker, som till exempel boende eller ekonomiska frågor.
Om du avser att bo i Finland i över tre månader, ska du ansöka om Registrering av uppehållsrätten för EU-medborgare hos Migrationsverket.
Du behöver inget mopedkort om du har fyllt 15 år före den 1 januari 2000.
Du kan boka en tid i förväg på Ajovarmas webbplats.
Du kan be om information om undervisning i finska och svenska för invandrare hos utlänningsbyrån.
Information om statsborgen för bostadslånfinska _ svenska _ engelska
Personer under 18 år och gravida har rätt att få alla de hälsovårdstjänster som övriga helsingforsare får.
Verksamhetsstället i centrum
På telefonen ger den jourhavande överinspektören råd om hur du kan utreda saken och kommer överens om eventuella fortsatta åtgärder för att föra saken vidare.
Att häva hyresavtalet omedelbart om det är skadligt för hälsan att bo i bostaden.
På ungdomsgårdarna har ungdomarna kostnadsfritt tillgång till ett mångsidigt urval av hobbyredskap, så utbudet av aktiviteter är stort.
Familjebandet mellan föräldern och barnet måste bevisas till exempel med en födelseattest med föräldrarnas namn.
Grundläggande utbildning för unga invandrare
FPA:s stöd är till exempel
Uppvärmning
Mer information finns på InfoFinlands sida Stöd till gravida.
Tågtidtabellerfinska _ svenska _ engelska _ ryska
linkkiSocial- och hälsovårdsministeriet:
linkkiStudentexamensnämnden:
Magistraterna (maistraatti) är lokala statliga förvaltningsmyndigheter.
Om du får lönen utbetalad i kontanter, ska du ge din arbetsgivare ett skriftligt intyg om löneutbetalningen.
MoniNet, som i Rovaniemi upprätthålls av Rovalan Setlementti ry, är ett center för mångkulturell information och verksamhet.
Du kan också söka ersättning från FPA i efterhand.
Om du ska arbeta i ett EU-/EES-land omfattas du av den sociala tryggheten i arbetslandet under den tid då du arbetar i landet, även om arbetet pågår mindre än sex månader.
Huruvida du beviljas uppehållstillstånd beror på hur starka och nära släktband du har till Finland.
Läs mer på InfoFinlands sida Företagsformer.
Frivilligarbete är inte samma sak som arbete eller praktik.
År 1765 erhöll staden stapelrättigheter, dvs. rätt till fri utrikeshandel, främst tack vare den aktiva kyrkoherden och lantdagsmannen Anders Chydenius.
Du kan söka till Finnish for Foreigners-kurserna via öppna universitetet.
Om det måste göras förändringsarbeten eller installeras fasta hjälpmedel i din bostad kan du få ersättning för detta av din hemkommun.
Vad bör jag göra?
Ni kan även välja att ta ett helt nytt efternamn som ert gemensamma namn.
Problem i äktenskap och parförhållande
Undervisningen kan bestå av närundervisning, distansundervisning, webbundervisning och självständiga studier.
Om du behöver särskilt stöd i de yrkesinriktade studierna t.ex. på grund av handikapp eller inlärningssvårigheter ska du ansöka till utbildningen via ansökan till specialundervisning.
Båda pensionssystemen omfattar ålderspension och invalidpension.
Vissa personer, till exempel äldre eller personer med funktionsnedsättning, har svårt att klara av de dagliga sysslorna utan hjälp.
Stöd och verksamhet för rörelsehindradefinska
hälso- och välbefinnandeområden
linkkiFinansbranschens Centralförbund:
Om du har studerat vid öppna universitetet och söker till universitetet ansöker du via separat ansökan (erillinen haku).
Om du har barn under 13 år och överväger att skilja dig, ta kontakt med familjerådgivningen (perheneuvola).
Helsingfors stad ordnar tjänster för personer med funktionsnedsättning, till exempel hjälpmedel, färdtjänst och dagverksamhet.
Boka en tid vid tjänstestället och ta med dig den ifyllda ansökningen, bilagorna och en identitetshandling.
försäkring
Småbarnspedagogik är avsedd för barn under skolåldern.
Arbetsgivaren betalar skatterna direkt från din lön.
linkkiHOAS:
Skilsmässa kan sökas av den ena eller av båda makarna tillsammans.
Ett innehavarkort (haltijakohtainen kortti) kan användas av flera personer.
Oftast söker man separat till dessa klasser.
Hur ordnas umgängetfinska
Checklista för den som ska färdas på isen:
Om en av makarna ensam ansöker om skilsmässa, börjar betänketiden från den dag då ansökan delges den andra makan.
Om du är medborgare i ett land utanför EU, måste du ansöka om uppehållstillstånd i Finland.
Hur beräknas skatteprocenten?finska _ svenska
Miljöministeriet linkkiMiljöministeriet:
Fritidsverksamhet för seniorer
Migrationsverket beslutar baserat på din berättelse om du beviljas asyl i Finland.
De stödjer sitt barns inlärning.
Också många privata företag erbjuder idrottshobbyer för barn.
Garantipensionen tryggar ett existensminimum för pensionärer.
Designmuseetfinska _ svenska _ engelska
äktenskapsintyg
Köp och sälj använda produkter.
Namnet på Finlands äldsta stad, Åbo (Turku), betyder handelsplats.
Ett brev som tillhör en annan person får inte läsas och en annan persons telefonsamtal får inte avlyssnas.
Om barnet eller den unga har flyttat till Finland nyligen, kan hen få förberedande undervisning före den grundläggande utbildningen.
linkkiSkattemyndigheten:
Diskrimineringslagen förbjuder diskriminering på grund av ålder, ursprung, nationalitet, språk, religion, övertygelse, åsikt, politisk verksamhet, fackföreningsverksamhet, familjeförhållanden, hälsotillstånd, funktionsnedsättning, sexuell läggning eller någon annan omständighet som gäller den enskilde som person.
Plötsliga krissituationer kan till exempel vara en allvarlig olycka, att en närstående avlider eller att du blir offer för våld.
Försörjningsförutsättning för make/maka/sambo/partner till en flykting
Alla familjemedlemmar kan inte få uppehållstillstånd.
Medborgare i EU- och EES-länderna kan anmäla sig som arbetslösa på nätet i TE-byråns ”Mina e-tjänster”.
På InfoFinlands sida Boende hittar du mer information om hur du söker bostad och andra frågor i anslutning till boende.
Kom ihåg att anmäla dig också direkt efter studier, arbetskraftsutbildning eller en period med sysselsättningsstöd.
Kvotflyktingarna väljs bland de personer som UNHCR föreslår till Finland.
Arbetstagare eller företagare
Rättshjälp till flyktingarfinska _ svenska _ engelska
Registrering som invånare
Stöd för hemvård av barnfinska _ svenska
på finska, tfn 029 502 4880
InfoFinland
Läs mer på InfoFinlands sida Ambassader i Finland.
Skatt som betalas direkt från lönen, är förskottsskatt (ennakonpidätys).
Du behöver också en finländsk personbeteckning.
Också barnet för vilket man söker underhållsstöd ska bo i Finland.
Finland tar som kvotflyktingar emot personer som har flyktingstatus enligt Förenta nationernas flyktingorganisation UNHCR.
avgångsbetyg från gymnasiet med ett godkänt vitsord i finska eller svenska som modersmål eller som andra språk
Föreningen för mental hälsa i Finland (Suomen Mielenterveysseura) har en kristelefon som ger samtalshjälp för människor i en krissituation.
Operationen görs på sjukhus och återhämtningen tar vanligtvis 1–2 dagar.
En inledande kartläggning och integrationsplan utarbetas för dig i arbets- och näringsbyrån. Om du kommit till
Stadens tjänster för arbetslösa
Kontaktuppgifter till tingsrättfinska _ svenska _ engelska
legaliserat äktenskapsintyg (om du är gift)
Man behöver inte be om tillstånd från till exempel släktingar.
Information om rättshjälpfinska _ svenska _ engelska
Äktenskap som ingåtts utomlands
Om du studerar utomlands och vill komma till Finland för arbetspraktik behöver du ett uppehållstillstånd på grund av praktik.
Öppettider: mån–fre kl. 9.00–16.00
Du kan meddela om avdrag, när du beställer ett nytt skattekort.
Om saken inte kan lösas på arbetsplatsen ska du kontakta arbetarskyddet vid Regionförvaltningsverket i Västra och Inre Finland.
Språkkaféerna är avgiftsfria.
Öppet alla dagar dygnet runt.
Länder där en annan Schengenstat representerar Finlandfinska _ svenska _ engelska
Tfn 029 56 60123 mån–fre kl. 8–16.15
På arbetsplatsen representeras fackförbundet och de anställda som är medlemmar i det av förtroendemannen.
Du kan också köpa ett prepaid-abonnemang.
Familjerådgivningen/familjecentret
Äktenskapsförordet skickas till magistraten för registrering.
Det är ofta svårt att uppskatta rätt belopp.
linkkiSanta Sport :
Vissa daghem och familjedagvårdare har öppet dygnet runt med anledning av föräldrarnas arbete eller studier.
Tfn: (09) 8392 4202
Vissa gymnasier är specialgymnasier.
Utländska beskickningar i Finland
Du hittar kontaktuppgifterna till Brottsofferjouren på webbplatsen.
Du kan fråga mer om kartläggningen och integrationsplanen vid utlänningsbyrån eller TE-byrån.
Vid läroanstalterna börjar kurserna vanligtvis i augusti eller september och i januari.
Barnfilmerna är ett undantag. De kan vara dubbade till finska även om filmens originalspråk är något annat.
Finland för en längre tid än för en kort semesterresa, ska du också anmäla detta till FPA (Kela) Om du omfattas av den sociala tryggheten i Finland och flyttar utomlands för högst ett år, bibehålls din rätt till den sociala tryggheten i Finland vanligen under din vistelse utomlands.
På webbplatsen för Finlands översättar- och tolkförbund finns en sökmotor med vilken du kan söka en tolk eller en översättare.
Folkhögskolan Työväen Akatemia tillhandahåller undervisning inom många akademiska discipliner samt träning för dem som vill läsa på universitet.
Lagen angående vårdnad om barn och umgängesrättfinska _ svenska _ engelska
Du har rätt till gottgörelse till exempel då varan som du köpt har fel som inte du har orsakat.
Rusmedelsbruk
personlig hjälp och dagverksamhet
Förfrågningar om bostadsrättsavgifter och bruksvederlag samt om lediga bostäder eller bostäder som kommer att bli lediga ställs direkt till ägaren.
Efter Nöteborgsfreden 1323 hörde största delen av det finska territoriet till Sverige.
Olika konstarter är musik, bildkonst, dans, teater och cirkuskonst.
Jämlikhet (yhdenvertaisuus) betyder att alla människor är likvärdiga oberoende av kön, ålder, etnisk eller nationell härkomst, nationalitet, språk, religion och övertygelse, åsikt, handikapp, hälsotillstånd, sexuell läggning eller någon annan orsak som gäller hans eller hennes person.
Du ska skaffa dig det europeiska sjukvårdskortet i det land där du har din sjukförsäkring.
Öppettider: mån–fre kl. 9.00–16.00
Inflyttningen till Esbo blev livligare från och med 1940-talet.
Övningar och kurser på internet
Information om att bo i delägarbostadfinska _ svenska _ engelska
Om du har ekonomiska problem kan du fråga om råd hos kommunens socialarbetare.
religion,
Barnatillsyningsmännenfinska _ svenska _ engelska
Hyrorna för Helsingfors stads hyresbostäder är lägre än de för privata hyresbostäder.
får utkomststöd eller
Barnrådgivningsbyråerna (lastenneuvola) och familjerådgivningsbyråerna (perheneuvola) ger råd i frågor som rör barns hälsa, uppväxt och utveckling.
Kelviå tandklinik
linkkiUtvecklingsstördas intressebevakningsorganisation:
Styrelsen ska bestå av minst ordföranden och två medlemmar.
Hemvård
Barnskyddslag
Tfn 029 56 60120
Studenterna tar på sig sina vita studentmössor.
Tjänster för småbarnspedagogik
Bland annat på internet och i dagstidningar finns det annonser för bostäder som är till salu.
Faderskapsledigheten är den del av föräldraledigheten som är avsedd att tas ut av fadern.
Hindersprövningen görs på magistraten (maistraatti).
InfoFinland är en webbtjänst på 12 språk där alla språkversioner är identiska.
Om du röstar på valdagen, kan du rösta endast på det ställe som anges på kortet.
Kipinä
familjeförhållanden
Läkemedel
Båda föräldrarna registreras som barnets vårdnadshavare.
Läs mer om ämnet på InfoFinlands sidor Stöd till gravida och Stöd efter barnets födelse.
Ett barn som har ett annat modersmål än finska eller svenska lär sig finska eller svenska som främmande språk.
Läs mer: Finska och svenska språket.
På Grankulla stadsbibliotek kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
Dessutom ska den ifrågavarande kommunen vara din hemkommun den 51:a dagen före valdagen.
Ansökan ska lämnas in fyra månader innan du behöver plats inom småbarnspedagogiken.
Läs på FPA:s webbsidor när familjeförmåner betalas ut till utlandet.
När du behöver hjälp av polisen i en nödsituation, ring det allmänna nödnumret 112.
Skilsmässa och uppehållstillstånd
Endast en läkare får utföra operationen.
Presidentkandidater kan nomineras av
Kommunerna har självstyre, vilket betyder att de själva kan besluta om ärenden i kommunen.
Bussbiljetterfinska _ svenska _ engelska
På studiepenningens belopp inverkar bland annat stödmottagarens ålder, om hen bor i sitt eget hem eller hos en förälder, on hen är gift och om hen har minderåriga barn. Kontrollera storleken på din studiepenning på FPA:s webbplats eller vid en FPA-byrå.
Hjälp och rådgivning
Vanligtvis kan du få handikappbidrag när du har bott tre år i Finland.
Finland har alltid varit en nordlig och liten plats mellan öst och väst.
Information om hyresboendefinska _ svenska _ engelska
På InfoFinlands sida Problem i äktenskap och parförhållande finns uppgifter om vart du kan vända dig för att få hjälp vid problem i parförhållandet.
Dagvård och förskoleundervisning
Säsongsarbetet kan pågå högst nio månader.
När ett barn föds, får barnet finskt medborgarskap om
Det innebär att du måste flytta ut ur bostaden och betala de obetalda hyrorna.
Finland ett självständigt land och den 6 december firas än idag som Finlands självständighetsdag.
Tandvård
Du kan få handledning i företagande eller företagarutbildning.
I InfoFinland finns information om tjänsterna i många kommuner.
Uppehållstillstånd för säsongsarbete
Yrkeshögskolafinska _ engelska
Om det inte finns någon uppgift om ditt civilstånd i Finlands befolkningsdatasystem, ska du lämna in ett ämbetsbevis (siviilisäätytodistus) från myndigheten i ditt hemland till magistraten.
En del av kurserna är avsedda för personer som vill grunda ett företag, och en del för dem som redan har ett eget företag.
När bodelningen inleds ska man utreda hur mycket egendom och skulder vardera maka har.
Nybörjarkurs i finska, Easyfinnishfinska
Kontaktpunkt för gränsöverskridande hälso- och sjukvårdfinska _ svenska _ engelska
Brottsutredning
På 1930-talet var många högersinnade och högerextrema rörelser populära i Finland liksom i det övriga Europa.
Delas egendomen jämnt eller inte?
Uppehållstillstånd för säsongsarbete
Läs mer på InfoFinlands sida Hemkommun i Finland.
Många organisationer erbjuder fritidsverksamhet och kamratstöd till personer i alla åldrar.
Ett par kan välja om de vill leva tillsammans i ett samboförhållande eller i ett äktenskap.
Läs mer: Museer.
prövotidens längd
Meritförteckning eller CV
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
Grannmedling innebär att grannarna diskuterar och en utomstående medlare leder samtalet.
Den förberedande undervisningen pågår vanligtvis i ett år.
I vissa fall får du en tolk genom myndigheten om du meddelar behovet av tolkning i förväg.
I Finland är det ofta svårt att hitta arbete om man inte kan finska eller svenska.
Tfn (09) 310 466 28
Om ditt företag har förutsättningarna för en lönsam verksamhet men du inte har tillräckligt mycket pengar eller säkerheter för att få ett banklån, ska du fråga om du kan få ett lån eller borgen hos Finnvera.
Rådgivning för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
Till att börja med görs en skriftlig skilsmässoansökan.
få finskt medborgarskap (18–22-åringar), om personen bott länge i Finland.
Ofta ska du betala en vattenavgift för bostaden.
Med läkaren eller psykologen kan du samtala konfidentiellt.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Permanent uppehållstillståndfinska _ svenska _ engelska
Vid problem kan du fråga råd hos arbetarskyddsfullmäktige eller förtroendemannen.
en syn- och hörselskada eller
För barn under skolåldern görs en tandläkarkontroll med ett par års mellanrum.
När du åker till sjukhuset ska du ta med dig tillräckligt varma kläder för barnet för hemresan.
Fyll i ansökningsblanketten i tjänsten Studieinfo.fi.
Du kan studera till exempel bland annat språk, estetiska ämnen, handarbete och kommunikation.
Äktenskapslagen finns i sin helhet på Finlex webbplats.
Orsaken till detta är arbetssäkerhets- och hygienföreskrifter som anknyter till arbetsuppgifterna.
Dagverksamhetfinska
Du kan registrera dig vid Helsingfors enhet vid magistraten i Nyland.
Registreringsintyget för den EU-medborgare, med vem du kommer till Finland
Information om allmänna insamlingsställen finns på adressen kierratys.info.
Ordna bokföringen
Också andra anhöriga till finska medborgare än en make/maka, en sambo, föräldrar till minderåriga barn eller minderåriga barn kan i vissa fall få uppehållstillstånd i Finland på grund av familjeband.
Invandrarenheten vid Helsingfors stads social- och hälsovårdstjänster hjälper invandrare bosatta i staden att integrera sig.
Regionförvaltningsverken sköter följande:
Kontaktuppgifter för förlossningsavdelningen:
Då pågår många evenemang på olika håll i Helsingfors.
Information om att söka arbete i Finland hittar du på InfoFinlands sida: Var hittar jag jobb?
Telefonnumret till Helsingfors Global Clinicin är 044 948 1698.
Kräv att arbetsgivaren betalar ut lönen.
Tfn 09 816 31300
Handbok för familjer med två kulturer (pdf, 4,74 Mt)finska _ engelska _ ryska _ franska _ spanska _ thai
I nödfall får du behandling även om du inte har en hemkommun i eller uppehållstillstånd till Finland.
Finland har haft svenskspråkig befolkning i över 800 år.
Det är obligatoriskt att registrera språket.
du är arbetslös arbetssökande
Min granne för oljud.
Drick kranvatten, det är gott och säkert i Finland.
Naturhuset är öppet för alla och ligger vid sidan av Bredvikens naturskyddsområde.
Åldersgränsen på ungdomsgårdarna varierar.
Samtidigt började man bygga Helsingfors innerstad i empirestil, vars byggnader inhyste storfurstendömets viktiga institutioner.
Eftermiddagsverksamhetfinska _ svenska
Dagvård fås på finska och på svenska.
Verksamheten utformas enligt ungdomarnas önskemål och de unga kan själva påverka innehållet i verksamheten.
Du får närmare anvisningar om hur du upprättar en affärsverksamhetsplan vid företagsrådgivningscentra.
I Esbo finns flera friluftsområden där man kan vandra i naturen.
Även en korrigerande operation är möjlig.
Vanda stads tjänster för invandrare (Vantaan maahanmuuttajapalvelut) ger dig information om integration, social- och hälsovårdstjänster och om stadens och olika organisationers tjänster.
Om du ska arbeta i Finland som specialist kan du även komma till Finland utan uppehållstillstånd.
Om Migrationsverket fattar ett negativt beslut på din asylansökan, har du rätt att arbeta under tiden då en eventuell överklagan behandlas.
Säkerhet och borgen för bostadslån
Dät är alltid bra att boka en tid i förväg på tjänstestället.
Det kostar i allmänhet att använda husbolagets bastu, tvättstuga och bilplatser.
Lediga jobbfinska _ svenska
Lapplands arbets- och näringsbyrå
Säkerheten är viktig till sjöss.
Guide till volontärarbetefinska _ engelska
Ni kan ta ett gemensamt efternamn om
Telefon: 09 816 31300
Ta kontakt med hjälpsystemet till offer för människohandel om du upplever att du blivit offer för utnyttjande.
Integrationsutbildningen är arbetskraftsutbildning och man söker till kurserna via Rovaniemi TE-byrå.
Om du behöver råd eller stöd för att hitta sysselsättning eller utbildning i finska språket, kontakta Helsingfors stads sysselsättningstjänster.
Du kan få låna olika hjälpmedel för att lättare kunna röra på dig, till exempel en käpp eller en rullator.
Arbetstagaren har rätt att på begäran få ett arbetsintyg av arbetsgivaren när anställningen upphör.
Av glaset tillverkas nya glasförpackningar.
Läkaren skriver vid behov en remiss till psykiatriska polikliniken (psykiatrian poliklinikka) eller en annan vårdenhet för psykisk hälsa.
Hjälp med rusmedelsberoendefinska _ engelska
Finsk personbeteckning
bostadens skick
Då tittar många finländare på självständighetsdagens mottagning med presidenten som värd på TV.
Om du inte fått ett brev om förskoleplats eller ansöker om förskoleplats under annan tid på året, ta kontakt med kontorstjänster för småbarnspedagogik per telefon på numret 040 806 5089.
Kommunen övervakar den privata småbarnspedagogiken.
Information om grundlagenfinska _ svenska _ engelska _ ryska
Handikappade personer
I Finland har många helgdagar rötterna i kristendomen.
Moninets webbplats
Anställningsrådgivning för invandrare
Sommarmånaderna i Finland är juni, juli och augusti.
Du kan fråga om råd vid socialbyrån (sosiaalitoimisto) eller rättshjälpsbyrån (oikeusaputoimisto) i din hemkommun.
hot, till exempel att hota med att skicka till hemlandet
Personen är skyldig att ersätta de skador som hen orsakat.
Undersökning av livmoderhalscancer görs på kvinnor i åldern 30–60 år vart femte år.
Hälsovårdstjänsterna i Esbo
I vissa situationer kan barnbidrag också betalas ut till utlandet, om du eller din make/maka omfattas av den sociala tryggheten i Finland.
I större städer kan det finnas apotek som har öppet till sent på kvällen.
Hobbygrupper finns både för nybörjare och mer avancerade.
Finland exporterade speciellt papper och andra produkter från skogsindustrin.
FPA:s ersättning kan ibland dras av direkt på det belopp som du betalar vid kassan.
Du måste ansöka om ett nytt uppehållstillstånd på grund av arbete innan ditt uppehållstillstånd för arbetssökande går ut.
Kontaktuppgifter:
Bostäder för ungdomar och studerande
Du hittar en lista över kurserna i finska på medborgarinstitutets webbplats.
Beslut om återkallande eller upphörande av uppehållsrätten fattas av Migrationsverket.
I Helsingfors finns även andra bibliotek, till exempel vid universiteten och högskolorna.
Yrkesutbildningen är mer praktiknära än gymnasieutbildningen.
Papper (paperi)
Beskickningen kan hjälpa dig om du har råkat ut för en olycka, blivit sjuk eller blivit utsatt för ett brott.
Dina familjemedlemmar kan inte få uppehållstillstånd i Finland på grund av familjeband.
På vissa orter har informationen om kurserna samlats på ett och samma ställe.
Alla kan få undervisning i den egna religionen eller i livsåskådningskunskap i skolan.
Fråga mer i din kommuns rådgivningstjänster.
Santa Sport Spa
I Karleby finns stadens daghem, gruppfamiljedaghem, familjedagvårdare samt barnklubbar.
Via rådgivningsbyråernas telefontjänst kan du boka tid på rådgivningsbyrån och fråga hälsovårdaren om råd beträffande graviditet och barns hälsa.
I juni och juli är det sommarlov.
Nybörjarkurs i finskafinska _ svenska _ engelska _ ryska _ kinesiska _ tyska
Bostadsansökan och bilagor
Rådgivningsbyråerfinska _ svenska _ engelska
Läs mer på InfoFinlands sida Hur kan man ansöka om finskt medborgarskap?
Handikappbidrag för barn under 16 år
Mer information om detta finns på InfoFinlands sida Arbetsintyg.
Information om uppehållstillstånd för studierfinska _ svenska _ engelska
Läs mer på InfoFinlands sida Yrkeshögskolor
Om det inte finns en förtroendeman på arbetsplatsen och du är medlem i facket, kontakta ditt fackförbund.
linkkiFinlands Röda Kors:
Ansökan är giltig i tre månader.
Var och en får fritt yttra sina åsikter i tal och skrift.
Information om området har sammanställts bl.a. i Hanhikivi-guiden som publicerats på finska, engelska, svenska och ryska.
Du ges möjlighet att lämna landet frivilligt.
Barnatillsyningsmannen bekräftar överenskommelsen om var barnen ska bo, vården av barnen, umgängesrätt och underhållsbidrag.
Du kan ge respons till beslutsfattarna och tjänstemännen till exempel via det elektroniska responssystemet.
Du har rätt till rehabilitering efter ett arbetsolycksfall.
läkare
Om du inte har rätt att använda de offentliga hälsotjänsterna kan du söka hjälp på en privat läkarstation.
Birkalands räddningsverk:
Om du misstänker att du har en könssjukdom, men har inga symtom, ska du kontakta din hälsostation.
Ansökan
Mer information om invaliditetspension och rehabilitering får du av FPA, din pensionsanstalt eller av företagshälsovården.
Handbok för handikappservicefinska _ svenska
Organisationen utför informations-, utbildnings och socialarbete i Finland.
På 1960-talet flyttade tusentals finländare till Sverige, eftersom det fanns mer jobb och betalades högre löner i Sverige än i Finland.
Information om mentalvårdstjänsternafinska _ svenska _ engelska
att tvinga någon till äktenskap.
Det finns även fritt finansierade delägarbostäder (vapaarahoitteinen osaomistusasunto).
Religioner i Finland
Skicka länken till ditt videoklipp och dina kontaktuppgifter till Infobanken till adressen infopankki@hel.fi.
Mer information om skolhälsovården finns på social- och hälsovårdsministeriets (Sosiaali- ja terveysministeriö) webbplats.
Kan hyresvärden i efterhand kräva att jag ersätter för brister som jag inte har orsakat?
Rådgivningarna för familjeplaneringfinska _ svenska
linkkiVanda vuxenutbildningsinstitut:
uppehållstillstånd
Ur ansökan bör även framgå hur länge och varför du studerar utomlands.
Läs mer om högskolor på InfoFinlands sida Universitet.
Information om den sociala tryggheten i Finland
linkkiArbets- och näringsministeriet:
Läs mer om beskattningen i Finland på InfoFinlands sida Beskattning.
I ett bostadsaktiebolag har du skyldighet att
Ofta ska man ange sitt löneanspråk i ansökningen.
Samtidigt kan ni också komma överens om underhållsbidraget, d.v.s. det ekonomiska stöd som den ena föräldern betalar för barnet.
Du kan inte få uppehållstillstånd för uppstartsföretagare i Finland utan ett positivt utlåtande från Business Finland.
Finland industrialiserades kunde finländarna sälja allt mer industriprodukter till utlandet.
Om du behöver icke-brådskande tandvård ska du ringa munhälsans centraliserade tidsbokningen.
Du ska också ingå en sysselsättnings- och integrationsplan med TE-byrån och delta i de tjänster och åtgärder som TE-byrån erbjuder åt dig.
Om du får andra sociala förmåner eller arbetsinkomster under arbetslösheten, är din grunddagpenning mindre.
På de flesta arbetsplatserna duar alla varandra oberoende av sin ställning.
Om du behöver sköta ett ärende med myndigheterna i ditt hemland ska du ta kontakt med ditt lands beskickning.
Om du har blivit utsatt för diskriminering kan du även ta kontakt med diskriminerings- och jämställdhetsnämnden (yhdenvertaisuus- ja tasa-arvolautakunta.
Du kan också studera på internet.
Om barnets mor och far inte är gifta och faderskapet inte erkänns, är barnet officiellt faderlöst.
Lämna inte tvättmaskinen eller diskmaskinen på när du går hemifrån.
Om du har ett FPA-kort (Kela-kortti) ska du ta det med när du besöker hälsovårdsstationen.
Filmfestivaler
Om du först planerar att flytta till Finland, läs mer på InfoFinlands sida Flytta till Finland.
utsökningen,
Sökning av hyresbostäderfinska
Tidtabeller, biljettpriser och linjekartor hittar du enklast på Matkahuoltos webbplats på finska, svenska och engelska.
ID-kortfinska _ svenska _ engelska
Branschspecifika myndigheter beslutar om rätten att utöva ett reglerat yrke eller använda en yrkesbeteckning.
Modern och fadern kan få flexibel eller partiell vårdpenning samtidigt om båda har förkortat sin arbetstid och tar hand om barnet under olika tider.
Ungefär 90 procent av finländarna har finska som modersmål.
Adress: Albertsgatan 25
Läs mer om tjänsterna för utvecklingsstörda på InfoFinlands sida Tjänster för handikappade.
Om du vill driva ett framgångsrikt företag i Finland, är det viktigt att du känner till den finländska företagskulturen.
Invånarlokalfinska _ engelska
Information om demokratin i Finlandfinska _ svenska _ engelska
Den utbetalas så länge som asylansökan behandlas.
Faderskapspenningen (Isyysraha) är avsedd för fadern då han tar hand om barnet.
Vanda är än idag en viktig trafikknutpunkt.
Du kan rösta i presidentval om du är finsk medborgare och fyller 18 år senast på valdagen.
Faderskapsledighet som tas ut efter föräldrapenningperioden kan delas upp i högst två perioder.
Ta reda på var den närmaste brandsläckaren finns.
du får finskt medborgarskap.
Flygplatsen har goda trafikförbindelser till exempel med bil, buss och tåg.
Lämna din ansökning till den beskickning eller visumcentral dit du ställer din ansökan.
Till de flesta fackförbund kan man också ansluta sig genom att fylla i en anslutningsblankett på fackets webbplats.
Barns och ungas problem
Hemvårdsstödets vårdpenning är lika stor för alla; beloppet påverkas inte av familjens inkomster.
I Finland utkommer många tidningar.
Läs mer om underhållsbidrag på InfoFinlands sida Familjer med en förälder.
Virussjukdomar, såsom herpes och kondylom, kan inte botas med läkemedel, men symtomen kan lindras.
Barnet eller den unga kan få förberedande undervisning före den grundläggande utbildningen under vilken han eller hon studerar finska (eller svenska) och vissa läroämnen.
Inom hälsovården har du rätt att bli betjänad på finska och svenska.
Vid universitetet kan du avlägga licentiatexamen (lisensiaatti) eller doktorsexamen (tohtori).
Du kan ansöka om barnbidrag från FPA antingen via FPA:s webbsidor eller med en pappersblankett.
Öppet programmeringsgränssnittfinska
Det finns vissa villkor för att få utkomstskydd för de arbetslösa och TE-byrån utreder om dessa villkor uppfylls i din situation.
Sök till en YH-examen i den gemensamma ansökan till högskolor på våren eller hösten Till många utbildningar är det möjligt att söka endast på våren.
JA: matavfall, även härsken mat, kaffesump, hushållspapper, skal från frukter etc.
Om du råkar ut för ett brott kan du be om hjälp vid *Brottsofferjouren.
Det betyder att det stadgas i lag vilken utbildning som krävs för dessa yrken.
Fundera på vilka som är dina kunder och vilka önskemål de har.
När du blir företagare, kan du få startpenning för att trygga försörjningen när företagsverksamheten precis har börjat.
I utrikespolitiken tvingades Finland under en lång tid balansera mellan Sovjetunionen och väst.
Vid musikinstitutet kan man musicera.
Barnets far är finsk medborgare, men modern är inte det och föräldrarna är gifta med varandra.
Arbetsgivaren har rätt att:
Kundgatan 3 A, 4:e våningen
Läs mer: Yrkesutbildning.
I Finland finns två pensionssystem som kompletterar varandra:
Om skilsmässa stadgas i äktenskapslagen.
behovet av bostad.
I Finland finns ett kommunalt bibliotek eller stadsbibliotek på alla orter.
mån–fre kl. 8.00–16.00 (för personligt möte måste du boka tid)
Avkomlingar till infödda finska medborgare
För att sköta ett juridiskt ärende kan man få ett rättsbiträde bekostat antingen helt eller delvis med statliga medel.
Till kommunens tjänster hör till exempel hälsovård och barndagvård.
Om du har ett körkort som utfärdats i ett land som är anslutet till Genève- eller Wien-konventionerna kan du köra med detta kort högst två år i Finland.
Flerspråkiga ordböckerfinska
inställt flyg på grund av strejk eller väderförhållanden,
Om videon väcker frågor hos dig kan du fråga mer av en expert.
Ditt sociala skydd när du flyttar utomlands
Mun- och tandhälsan påverkar hälsan i hela din kropps hälsa.
Arbetsdiskriminering är ett brott.
Det är möjligt att avlägga högskolestudier vid öppna universitet och öppna yrkeshögskolor.
du genomgått läkarundersökning före utgången av fjärde graviditetsmånaden
Konvaljvägen 21
fängelse och tortyr
internationellt skydd
Fackförbunden strävar efter att trygga sina medlemmars intressen och rättigheter, försöker förbättra lönerna och anställningsskyddet samt förbättra arbetslivets kvalitet.
du behöver startpenningen för din försörjning
Vad kan jag studera i yrkesinriktad arbetskraftsutbildning?
Finska på arbetsplatsen
Även i vanliga grundskolor kan det finnas några klasser där undervisningen sker på ett främmande språk.
Invånarparker och klubbar
När du söker hjälp hos en jurist, är det bra att säkerställa att juristen har sakkunskap i det område där du behöver hjälp.
I Finland tar hindersprövningen ungefär en vecka.
Information om studiestödetfinska _ svenska _ engelska
Tfn (09) 871 4043
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska
Ibland behövs sjukhusvård.
Efter grundskolan kan du studera på gymnasiet eller en yrkesläroanstalt.
Telefon: (06) 8287 580
De planerar sin verksamhet och sin ekonomi ett år fram i tiden.
Kontrollera alltid med hyresvärden vilka möbler som ingår.
Tfn (09) 622 4322.
Information om den sociala tryggheten i de nordiska ländernafinska _ svenska _ engelska _ norska
Staden underhåller cykelvägar, motionsrutter, joggingbanor, skidspår, badstränder, bollplaner och skridskobanor samt platser för närmotion.
Då stiger den månatliga avgiften eller också förlängs lånetiden.
Hälsostationerna har stängt kvällstid och under veckoslut.
Mentalvårdstjänsterfinska _ svenska
I Finland är det inte vanligt att visa sina känslor offentligt.
JA: lysrör, energibesparingslampor, kemikalier med ett varningsmärke på förpackningen
Religion
Jämställande av nivån på en högskolexamen
inte är gift eller i registrerat parförhållande sedan tidigare.
Avtala med din tjänsteleverantör om överföringen av din internetanslutning i god tid så att det inte blir ett avbrott i servicen.
Målet är att familjen meddelas om dagvårdsplatsen senast två veckor innan dagvården inleds.
linkkiDreamwearclub ry.:
Om du redan har haft ett uppehållstillstånd i Finland, men tillståndet inte förlängs, fattar Migrationsverket beslut om utvisning.
Mer information finns på Helsingfors vuxengymnasiums webbplats.
FPA:s pensioner utomlands
I Finland ordnas årligen högklassiga filmfestivaler, varav de bäst kända är Kärlek och anarki-festivalen, som ordnas varje höst i Helsingfors, och Sodankylä filmfestival som ordnas på sommaren.
Stöd till flyktingarfinska _ svenska _ engelska
I planen nedtecknas vilket kunnande du har förvärvat tidigare och fastställs vilka studier du ska avlägga.
Sjukvård
fre kl. 8–15.30
Bidrag och priserfinska _ svenska _ engelska
linkkiFCC, STTK och AKAVA:
Utlänningar ska enligt lag anmäla till registret samma uppgifter som finska medborgare om deras vistelse i Finland varar över ett år.
Om du flyttar till Finland för att bo här stadigvarande i ett år eller längre, ska du också registrera dig i magistraten på din hemort.
När du ska besöka tjänstestället, ta med dig din ifyllda ansökan, bilagorna och kopior på bilagor samt pass och passfoto.
Patientombudsmannenfinska _ svenska _ engelska _ ryska
Du kan ha rätt att få stöd från ditt eget hemland.
Du hittar mer information om den sociala tryggheten i Finland på FPA:s webbplats och på InfoFinlands sida Den sociala tryggheten i Finland.
Man får oftast en privat hyresbostad snabbare än en kommunal hyresbostad. Hyran för en privat bostad är ofta högre.
Det humanistiska och pedagogiska området
Barn till föräldrar i samboförhållande
Mer information om att köpa en egen bostad får du på banken eller hos fastighetsförmedlare.
Ditt anställningsavtal
Korso hälsostation, Fjällrävsstigen 6
Man kan anmäla sig till förskoleundervisningen antingen elektroniskt eller med en ansökningsblankett.
Rådgivningen ges på många olika språk.
Hälsovårdaren antecknar uppgifter om barnets hälsa och vaccinationer på kortet.
Arbetsgivaren kan utöver de lagstadgade försäkringarna även teckna olika frivilliga försäkringar åt sina anställda.
linkkiMuseiverket:
Om du inte har en hemkommun i Finland, räknas du som invånare i den kommun där du vistas.
Invandrarenhetens tjänster är till exempel vägledning, rådgivning och inledande kartläggning.
Du kan läsa mer om registrering av barnets födelse, faderskapserkännande och vårdnaden om barnet på InfoFinlands sida: När ett barn föds i Finland.
får kontakter till det finländska samhället.
Utöver dagsgymnasierna som är avsedda för ungdomar finns det tre vuxengymnasier (aikuislukio) i Helsingfors.
Öppet mån–fre kl. 8–16.15
Om du inte bor stadigvarande i Finland och blir utan bostad, ta då kontakt med ditt lands beskickning i Finland.
linkkiHumanistiska yrkeshögskolan:
Var även direkt i kontakt med TE-byrån om du önskar ändra en tidsbokning.
Den nuvarande regeringenfinska _ svenska _ engelska
Hjälp till offer för familjevåldfinska
Köpebrevet är ett kontrakt där t.ex. bostadens pris, bostadens storlek, bostadens skick och datumet då köparen får tillgång till bostaden finns inskrivet.
Kulturbranschen (musiker, inredningsarkitekt)
Anvisning om brottsanmälanfinska _ svenska _ engelska
Läs mer: Prövning av hinder mot äktenskap, Äktenskap
Om uppgifterna inte är korrekta, eller om det saknas något, komplettera och korrigera skattedeklarationen i webbtjänsten MinSkatt.
dina barns födelseattester.
Per post får du från EES-länderna beställa den mängd läkemedel som motsvarar högst tre månaders förbrukning.
Mentalvårdstjänsterfinska _ svenska _ engelska
Regionförvaltningsverket i Västra och Inre Finlandfinska _ svenska _ engelska
Vid institutet kan du avlägga enskilda kurser eller studera på någon av institutets studielinjer.
Du hittar bostäder till försäljning på sidor för bostadssökande på internet.
Inkassobyrån skickar dig genast ett betalningskrav.
Närmare information om hur man ansluter sig till avtalet ger InfoFinlands chefredaktör Eija Kyllönen-Saarnio, eija.kyllonen-saarnio(snabel-a)hel.fi, tfn 050 363 3285.
Arbetstagaren har rätt att få en lönespecifikation där det står vad lönen består av.
Apoteken har vanligen öppet från morgon till kväll.
Till småbarnspedagogiken hör mångsidig verksamhet, till exempel lekar, motion, utevistelse, musik, pyssel och utfärder.
För varje studerande utarbetas ett eget studieprogram.
Begravningsplatserfinska
Säsongsarbete är till exempel:
När du har fått ett läkarutlåtande eller en rehabiliteringsplan kan du ansöka om rehabilitering vid din arbetspensionsanstalt eller FPA.
Barn lär sig nya språk snabbt, även om det kan kännas svårt i början.
På magistraten utreder man även om det är möjligt att registrera en hemkommun i Finland för dig.
Utbildning för invandrarefinska _ engelska
Stationsbron i Esbo
Framför kravet skriftligt.
Vilka försäkringar måste jag ha?
Det närmaste förlossningssjukhuset är Jorv sjukhus i Esbo.
Under denna tid förlorar du inte rätten till invaliditetspension.
Om barnet har ett annat modersmål än finska eller svenska kan kommunen ordna undervisning i barnets eget modersmål.
linkkiInformationscentralen för teater i Finland:
religion.
På InfoFinlands sida Finska och svenska språket hittar du information om möjligheterna att studera finska eller svenska.
Att hälsa
Hurdant är det svenska språket?
Den vanligaste företagsformen är en enskild näringsidkare, vilket betyder att man driver företagsverksamhet utan ett skilt grundat företag.
Ett andelslag kan ha en eller fler medlemmar.
Om barnet har en hemkommun i Finland, kan du ansöka om Fpa-stöd för privat vård.
Berätta också hurdan bostad du letar efter.
I slotten ordnas också guidade rundvandringar där slottets historia och arkitektur presenteras.
Läs mer på InfoFinlands sida Hälsovårdstjänster i Finland och Hemkommun i Finland.
Om du upplever diskriminering på arbetsplatsen ska du först ta kontakt med din förman.
Barnatillsyningsmannenfinska _ svenska
Till HelMet-biblioteket hör även biblioteken i Esbo, Vanda och Grankulla.
Ring 112 till exempel i följande situationer:
Detta är ändå inte alltid fallet.
Tjänsten har öppet måndag till fredag kl. 9.00–16.00.
Bostäder för ungdomar och studerande
Om du har en betalningsanmärkning, får du inte nödvändigtvis en hyresbostad, ett banklån eller ett kreditkort.
Du behöver en hemkommun för att kunna använda kommunala tjänster, såsom hälso- och sjukvården eller dagvården.
I det ingår nästan alltid rätt att arbeta.
Ett efternamn som maken eller makan har fått från sitt tidigare äktenskap kan inte väljas som efternamn.
I Finland gör läkare inom de offentliga hälsovårdstjänsterna inga hembesök.
Information om förskoleundervisningenfinska _ svenska _ engelska
Om barnet är frånvarande från skolan till exempel på grund av sjukdom ska du meddela skolan om detta på morgonen via Wilma.
linkkiAndra ämbetsverk:
barn till syskon (till exempel morbror och systerdotter).
Sjukanfall och olyckor
Stöd för mångkulturella familjerfinska _ svenska _ engelska
Bibliotekets webbtjänstfinska _ svenska _ engelska
Din situation bedöms i sin helhet.
På apoteket kan du byta ut det läkemedel som föreskrivs på receptet mot ett annat, förmånligare läkemedel om det verksamma ämnet är detsamma i båda preparaten.
Rovaniemi stad/kulturtjänster linkkiRovaniemi stad/kulturtjänster:
linkkiDuo För bikulturella familjer:
FPA ger mer information om förtida ålderspension och tilläggsdagar till folkpension.
Av kartong görs exempelvis papprullar för hushållspapper.
Du får närmare uppgifter från tjänsten Studieinfo.fi.
När du blir sjuk ska du kontakta hälsostationen (terveysasema) på din ort.
Barnatillsyningsmannens tjänster hjälper föräldrarna att vid skilsmässa komma överens om avtal som är i barnets intresse.
du har fått tillfälligt skydd
Information om den sociala tryggheten i Finland för EU-medborgarefinska _ svenska _ engelska
Adress: Kaisaniemigatan 4 A, vån. 6
Om den ena maken inte förvärvsarbetar ska den förmögnare maken stå för kostnader för till exempel mat och kläder.
Vid Väestöliitto får du information om föräldraskap.
Utöver sport har ungdomar också tillgång till många konstaktiviteter, som till exempel bildkonst, musik eller teater.
Kontaktuppgifter till magistraten i Helsingfors:
Företagshälsovårdsläkaren avgör om du kan deltidsarbeta medan du är sjuk.
Vid val av invånare till stadens hyresbostäder prioriteras de sökande som har ett akut bostadsbehov.
Mer information om jourmottagningarna hittar du på Vanda stads webbplats om hälsovårdstjänster.
Tfn 029 564 4000
Information om besöksförbudfinska _ svenska _ engelska
Den unga själv eller föräldrarna kan också kontakta familjerådgivningen.
Du behöver inte ringa eller besöka TE-byrån om du inte uttryckligen ombes göra detta.
Mer information om att söka arbetslöshetsersättning hittar du på sidan Arbetslöshetsförsäkring.
Global Clinic anmäler inte kunderna till polisen eller andra myndigheter.
Öppna universitetet
På Esbo stads webbplats finns kontaktuppgifterna och telefonnumren till hälsostationerna.
På skattebyrån kan du till exempel få skattekort, ändra din skatteprocent eller fråga om sådant som rör beskattningen.
Delta och påverkafinska _ svenska
Det behöver du när du ansöker om moderskapsunderstöd (äitiysavustus) och moderskapspenning (äitiysraha) hos FPA (Kela).
Det innebär kortvarig (2–3 tim. per gång) vård av småbarn ute i en lekpark.
Att ansöka om medicinsk rehabiliteringfinska _ svenska _ engelska
Att grunda ett företag.
Exempelvis i Konst-Vionoja-centret presenteras konstnären Veikko Vionojas verk.
Parkering
Lämna inte mat på en het spis utan uppsikt.
I skolorna i Vanda ges hemspråksundervisning i flera olika språk.
I Finland flaggar man på bestämda dagar som är intagna i kalendern.
Sedan får du ett yrkesbevis som bevisar din yrkeskunnighet.
Österbottens tingsrätt Karleby kansli
Du kan kontakta rådgivningen om ditt barn har problem eller om ni har problem i familjen och du vill ha hjälp.
Fråga hos FPA om du har rätt till bostadsbidrag eller något annat understöd.
Efter föräldraledigheten kan antingen modern eller fadern ta ut en oavlönad vårdledighet för att ta hand om barnet tills barnet fyller tre år.
Före flytten till Finland
Fråga din arbetsgivare vad företagshälsovården på din arbetsplats omfattar.
Läs mer på InfoFinlands sida EU-medborgare.
Under samtalet ställs frågor om de händelser och orsaker som tvingade dig att lämna ditt hemland.
Om ni har barn och beslutar er för att skiljas ska ni boka en tid hos barnatillsyningsmannen (lastenvalvoja).
studier
Utvecklingsstördas intressebevakningsorganisationfinska _ engelska
Ansvarsområdena övervakar att de lagenliga arbetarskyddsföreskrifterna följs på arbetsplatserna.
Dessutom krävs det i allmänhet att ditt uppehållstillstånd är giltigt, om du är skyldig att ha ett uppehållstillstånd.
Det är bra att informera förlossningssjukhuset på förhand om omskärelsen så att det kan beaktas vid förlossningen.
Karlebynejdens Utveckling Abfinska _ svenska _ engelska
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
Biografer
Mer information om flytt, uppehållstillstånd och personuppgifter fås från bland annat magistraten, polisen och invandrarbyrån.
Du behöver inte ansöka separat om måltidsstödet.
Du kan söka färdtjänst hos en socialarbetare inom handikappservicen i din hemkommun.
Vid krismottagningen får du hjälp och stöd i svåra situationer.
När ett barn insjuknar
Hjälp för män för att sluta med våldsamt beteendefinska _ engelska
Företagshälsovården kan du besöka under arbetstid.
Du kan ta körkort i Finland när du har fyllt 18 år.
Invandrare ges rabatt på vissa kurser.
stöd avsedda för barnfamiljer.
Uppgifter som registreras är bland annat namn, födelsedatum, medborgarskap, familjeförhållanden och adress.
På InfoFinlands sida Var hittar jag jobb?
På skatteförvaltningens webbplats finns mycket information om beskattningen i Finland.
Den är avsedd för invandrare.
Regionförvaltningsverket i Västra och Inre Finland
Varifrån kan jag få hjälp vid konflikter med min granne?
I Finland ligger medeltemperaturen på vintern under noll Celsiusgrader och på sommaren över +10 Celsiusgrader.
Telefonnumret är (09) 310 44222
Fullmäktigeledamöterna representerar olika politiska grupper.
På InfoFinlands sida Var hittar jag jobb? får du information om hur du söker arbete i Finland.
Problem i arbetslivet
Läs mer på InfoFinlands sida Ekonomiskt stöd och under rubriken När du vårdar en närstående i hemmet på sidan Äldre människor.
Löneanspråk
Ring nödnumret 112 om det är fråga om en nödsituation.
Alla Esbobor får fritt fiska med metspö och pimpla.
Kontrollera villkoren för pensionärsrabatten på biljettkontoren.
Företagslagstiftningfinska
Olika kurser ordnas för både barn och vuxna.
Väestöliitto tillhandahåller rådgivning telefonledes och via e-post när du behöver samtalsstöd i frågor som rör barnuppfostran eller relationerna i familjen.
Du har rätt till nödinkvartering och mathjälp om du inte har pengar till mat eller någonstans att övernatta.
En flykting är en person med flyktingstatus.
Ta kontakt direkt med den organisation där du vill arbeta som frivillig.
Förskoleundervisningen är avsedd för sexåringar och den ges vid daghem.
I A-klinikstiftelsens webbtjänst Päihdelinkki får du information om missbruk och beroende.
Yrkeshögskolorfinska _ svenska _ engelska
Information om rådgivningsbyråernas tjänsterfinska _ svenska _ engelska _ ryska
För att kunna arbeta i Finland behöver du vanligen antingen ett uppehållstillstånd för arbetstagare eller någon annan typ av uppehållstillstånd för förvärvsarbete.
Rådgivningen är avgiftsbelagd.
FPA:s ersättning kan ibland dras av direkt på det belopp som du betalar vid kassan.
Tillstånd för säsongsarbetefinska _ svenska _ engelska
I Karleby finns biografen Bio Rex, vars två salar använder digital- och 3D-teknik.
Förutom finska och svenska talas även andra inhemska språk i Finland.
Om du kommer från ett land som inte är ett EU-land, ett EES-land eller Schweiz till Finland för att studera behöver du vanligtvis ha en täckande sjukförsäkring i ditt hemland för att få uppehållstillstånd i Finland.
Kurdiska
Också punktlighet är viktigt för finländarna.
Vanda stad ordnar även klubbar (kerho) för 2,5–5-åriga barn som vårdas i hemmet.
Alla personer som har en adress i Finland kan få ett bibliotekskort.
Ellfolkgatan 5
I de flesta gymnasieskolorna är undervisningsspråket finska eller svenska.
Även medborgare i EU-länder och nordiska länder och deras familjemedlemmar har rätt att arbeta och studera.
Detta förutsätter att din arbetstid och lön uppfyller minimikraven.
Du måste hitta en arbetsgivare som vill anställa dig.
För annat fiske behöver du ett avgiftsbelagt tillstånd.
linkkiTullen:
TE-byrån ordnar
Begär bekräftande av avtalet hos barnatillsyningsmannen i din hemkommun.
Företagare i Finland
I Vanda finns också privata tandläkare.
Nyheter på ryskaryska
Asukastila Myyrinki
Stadsfullmäktiges sammanträden på Internetfinska _ svenska
Din kultur, ditt språk och din religion kan fortfarande utgöra en viktig del av ditt liv också i Finland.
Friluftsliv i skärgårdenfinska _ svenska _ engelska
Läs mer på InfoFinlands sida Företagsrådgivning.
Kommunernas verksamhetfinska _ svenska
Det är vanligt att man äter två varma måltider om dagen, lunch och middag.
Hälsa
linkkiArbetsministeriet:
Medarbetarna pratar finska, svenska och engelska.
Lapplands yrkeshögskolafinska _ engelska
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
Stöd för studierna och tionde klassen
Stadin asunnotfinska _ svenska _ engelska
Gymnasiet tar 2–4 år, beroende på den studerande.
Nödfall
Kontaktuppgifter till socialarbetarefinska _ svenska _ engelska
Ambassader och konsulat är statliga beskickningar i en annan stat.
Du kan ta ut vårdledighet om du har befunnit dig i samma arbetsgivares tjänst under minst 6 månader under det senaste året.
Där får du även en mall för affärsverksamhetsplanen och andra dokumentmallar.
Om du vill flytta ut ur bostaden måste du göra en avträdelseanmälan (luopumisilmoitus) till husets ägare.
I evenemangskalendrarna hittar du information om filmfestivaler i Helsingfors.
alla dina arbetsintyg och studiebetyg
Det är inte tillåtet att beträda folks gårdar utan lov.
Ansökan om uppehållstillstånd
Öppettider och kontaktuppgifterfinska
Jag talar bara lite finska.
Du lär dig språket bäst om du vågar använda det.
Förarutbildning kan du få i en bilskola.
Läs mer om tjänsterna för handikappade och om att ansöka dem på InfoFinlands sida Tjänster för handikappade.
Det kan också vara en hälsorisk att köpa läkemedel i en olaglig webbutik.
Läs mer: Teater och film.
Sjukpensionfinska _ svenska _ engelska
Finländare använder inte skor inomhus.
Såväl män som kvinnor och barn kan vara offer till människohandel.
Tfn (09) 272 2775 och 040 501 3199.
Skolbarns hälsa
Historia
Jag förstår inte, kan du upprepa?
Sverige och Ryssland stred under denna tid ett flertal gånger om vem som skulle vara makthavaren över Finland.
Du kan också besöka FPA:s kontor.
Om du har avlagt examen i något annat land kan du behöva beslut om erkännande av examen för att kunna arbeta eller studera i Finland.
barnets mor är finsk medborgare,
Uppskattningen baseras på beloppet av de beskattningsbara inkomsterna året innan.
Den gamla huvudstaden Åbo förstörs i en brand och Helsingfors får en allt viktigare ställning
Om du har fyllt 58 år innan du blev arbetslös, kan du få grunddagpenning i mindre än 500 dagar.
Om du har fyllt 70 år och Vanda är din hemkommun kan du kostnadsfritt använda Vanda stads simhallar och gym. Du kommer gratis in till idrottsanläggningarna om du har ett Sportkort (Sporttikortti).
Adress: Bangårdsvägen 7 (ingång via Loktorget)
Invandrare får hjälp med jobbsökningen vid Lapplands arbets- och näringsbyrå (TE-byrån).
Du ska vistas lagligt i det land där du ansöker om visum.
1968 Den finländska grundskoleinstitutionen inrättas
Förtroendemannen agerar som förhandlare, medlare och informationsförmedlare mellan arbetsgivaren och anställda.
Stödboende
Om du är intresserad av en bostad ska du kontakta något av de företag som tillhandahåller bostadsrättsbostäder:
Försörjningsförutsättning för make/maka till en utländsk medborgare
mottagningstjänster för invandrare
I ett kombinerat efternamn syns båda efternamnen, till exempel Virtanen-Smith.
Information om Finland
Äktenskap ingås genom vigsel.
Du får ett elavtal genom att ringa upp elbolaget och meddela ditt namn och din nya adress.
Läs mer på webbplatsen för linkkiFörbundet för mödra- och skyddshem:
Om man vill fortsätta studierna därefter och avlägga högre yrkeshögskoleexamen, måste man först skaffa sig tre år av arbetserfarenhet från samma område som examen.
Telefon: 040 1817 400
Yrkesutbildning
Seniorbostäderfinska _ svenska
Då får du ett graviditetsintyg av läkaren eller från rådgivningen.
Du kan anmäla dig antingen via nättjänsten eller personligen hos TE-byrån.
Du kan även gå till Vanda skyddshem eller huvudstadsregionens skyddshem.
Uppehållstillstånd för arbetstagarefinska _ svenska _ engelska
I lagstiftningen och kollektivavtalet fastställs till exempel minimilöner, arbetstider, semestrar, lön för sjukdomstid och uppsägningsvillkor.
arbetsförmedling
Vilka tillstånd behöver du?(pdf, 384 kt)finska _ engelska
I takt med industrialiseringen började flyttrörelsen från landsbygden till städerna.
Akutmottagningen
Du hittar grundläggande information om att starta ett företag i Finland på dessa sidor i InfoFinland.
Barnavård och hemhjälpfinska
Den person som får flest röster vid andra valomgången väljs till president.
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
I Vanda finns många politiska föreningar, invandrarföreningar och andra föreningar via vilka du också kan påverka beslutsfattandet.
När anställningen upphör har arbetstagaren rätt att få semesterersättning för de dagar som han eller hon inte har fått semester eller semesterersättning för vid tidpunkten för anställningens upphörande.
I beskattningen kan du göra avdrag (vähennykset), som minskar beskattningen.
Telefon: (06) 8264355.
På Utbildningsstyrelsens webbplats finns en förteckning över de reglerade yrkena och de ansvariga myndigheterna.
Om du behöver en tolk, skaffar Migrationsverket tolken.
För företagare är självrisktiden oftast dagen för insjuknandet och följande tre vardagar.
Serviceboendet omfattar både bostaden och tjänsterna som anknyter till boendet.
Läs mer: Vård av barnet
Sök lediga jobb på jobbförmedlingssidor på internet, i tidningar eller på sociala medier (till exempel Facebook och LinkedIn).
vigselbevis
du avlägger en kompletterande utbildning eller en specialutbildning som hör till din examen.
Arbetstagarnas inskolning och säkerhet
Kvinnor och män kan själva besluta om vem de gifter sig med.
FPA ger rådgivning på telefon även på ryska och arabiska.
Hyresbostäderfinska
Samjourens adress:
Arbetsavtalet kan vara tidsbundet om det finns en välgrundad orsak till detta.
Gymnasierfinska _ svenska _ engelska
Var får jag hjälp?
Ett barn kan födas utom äktenskapet eller också är dess föräldrar skilda.
Om ditt barn har hemkommun (kotikunta) i Finland har han eller hon rätt att utnyttja de offentliga hälsovårdstjänsterna.
Ett exempel på diskriminering är om du inte får betjäning på grund av ditt etniska ursprung eller om man vid en arbetsintervju kräver att du ska behärska finska språket fullständigt trots att det inte är nödvändigt i arbetet.
Namnen kan även skrivas isär, utan bindestreck.
Däremot kan man dela upp föräldraledigheten så att modern eller fadern stannar hemma växelvis för att ta hand om barnet.
Information om stöd till barnfamiljerfinska _ svenska _ engelska
Läs mer på InfoFinlands sida EU-medborgare.
Inhemska minoritetsspråk
Fråga mer om hobbymöjligheterna, tidtabellerna och priserna direkt hos arrangören.
Takorganisation för somaliska föreningarfinska _ engelska _ somaliska
Tjänsterna är avsedda för invandrare i Helsingfors som fyllt 17 år och har uppehållstillstånd.
Till exempel ett stambyte kan kosta bostadsägaren många tiotusentals euro.
Om du behöver en gynekologisk undersökning, ta kontakt med hälsostationen.
Elektronisk tidsbokningfinska _ svenska _ engelska
Avfallshantering i bostaden
Det är viktigt att komma ihåg att man inte får ge tobak eller alkohol till barn under 18 år.
Invandrareleverna bedöms som regel enligt grundskolans allmänna bedömningsgrunder med beaktande av elevens utgångsläge.
Krishjälpfinska _ svenska _ engelska
Puh. 040 126 7513
I Esbo finns simhallar, flera idrottshallar, idrottsplaner och andra idrottsplatser för olika idrottsgrenar.
Mina e-tjänsterfinska _ svenska
På bastulaven sitter man oftast på ett litet sittunderlag.
Om du behöver information om tillståndsärenden som sköts av polisen, fordonsföreskrifter eller hur undersökningen i ett brott som skett tidigare framskrider ska du ringa polisens egna nummer under tjänstetid.
intyg på yrkesinriktad grundexamen som du har avlagt på finska eller svenska
Äktenskapsförordet kan upprättas före eller under äktenskapet.
Att ansöka om sjukdagpenningfinska _ svenska _ engelska
– Du kan även lyfta fram dina intressen.
tfn 020 741 4732
Ytterligare information om yrkesutbildningfinska _ svenska
Vegetarism har blivit allt populärare.
Diskussionsgrupp på finskafinska
Om ni behöver hjälp med att komma överens om sådant som rör barnen kan ni ansöka om medling i familjeärenden.
Utbildning – Lista dina examina i kronologisk ordning, den senaste först.
linkkiYrkesläroanstalten Varia i Vanda:
Du får själv bestämma vilket trossamfund ditt barn ska höra till.
Gruppfamiljedaghemfinska _ svenska
Om du misstänker att du är offer för människohandel, kontakta systemet för hjälp till människohandelns offer (Ihmiskaupan uhrien auttamisjärjestelmä).
I Finland kan du studera på finska, svenska och ibland även på engelska.
Om du har rätt till hemvårdsstöd kan du ansöka om det vid FPA.
Om du har blivit utsatt för ett brott, kan du få hjälp och råd vid Brottsofferjouren.
Beslut i viktiga kommunala ärenden fattas av kommunfullmäktige (kunnanvaltuusto).
Du kan också få handledning i datoranvändningen och på vissa bibliotek ordnas finska språkcaféer.
Uppgift till myndigheterna i det egna landet (utländska medborgare)
Kurser vid folkhögskolor för invandrarefinska
För att få ett uppehållstillstånd för studerande, ska du kunna visa att din ekonomiska situation ger dig möjlighet att leva i Finland.
Du behöver personbeteckningen till exempel för din arbetsgivare eller läroanstalt.
Den förberedande utbildningen är avsedd för ungdomar och vuxna som är intresserade av yrkesutbildning och vill förbättra sina kunskaper i finska.
Tfn (09) 8195 5360
Stödtjänster för handikappadefinska _ svenska _ engelska
Begravningsbyråerfinska _ svenska _ engelska
Föräldrapenning till modern eller fadernfinska _ svenska _ engelska
Webbsidorfinska _ svenska _ engelska
Per telefon får du betjäning på finska, svenska och engelska.
Eventuella arbetsintyg (om du inte ska avlägga examen eller är en utbytesstudent)
Hyrarbetsguidefinska _ svenska _ engelska
Det kan vara svårt att hitta en bostad eftersom efterfrågan på bostäder är större än utbudet speciellt i större städer.
Företagare kan ordna sin egen företagshälsovård om de vill.
Kommunerna tillhandahåller tandvård vid hälsostationer (terveysasema) och tandkliniker (hammashoitola).
Tfn: 029 512 000
Läs mer Registrering som invånare
Du kan ansöka om tillståndet på internet i tjänsten Enter Finland.
Om du vill grunda ett eget företag, kan du få hjälp vid FöretagsEsbo.
Det finns också särskilda Erasmus Mundus-magisterprogram som har ett eget stipendiesystem.
Läs mer på InfoFinlands sida Kan jag förlora mitt uppehållstillstånd?
Allmän språkexamen
En del rutter är belysta.
Öppettider: varje dag kl. 17.00–10.00
Det kan vara svårt att komma in dit.
Skicka in en ansökan om namnändring till magistraten.
Telefonrådgivning av en jurist 0800 161 177
Barnets födelseattest om du har vårdnaden om ett barn
Anhållan om prövning av hinder mot äktenskapfinska _ svenska
Infomöten ordnas på finska, engelska, ryska, arabiska och estniska.
TE-byrån (TE-toimisto) hjälper dig att söka arbete.
I Finland finns också ett eget teckenspråk.
fostran
När du besöker magistraten, ta med dig minst följande handlingar:
Också en person kan vara ett hushåll.
Du hittar kontaktuppgifterna på diskrimineringsombudsmannens webbplats.
Tammerfors
Man kan ansöka om att omfattas av det finska socialskyddet av FPA då uppehållstillstånd har beviljats.
Nya barnsjukhuset (Uusi lastensairaala)
I Finland är enligt lag personer under 18 år barn.
Du får börja arbeta först när du har fått ett uppehållstillstånd.
Helsingfors och Sveaborg erövrades av ryssarna 1808 och under kriget brann staden.
Skatter betalas på de inkomster som företagaren eller företaget har kvar när alla kostnader för företagsverksamheten har dragits av försäljningen.
att tvinga någon till arbete, för vilket man betalar för lite eller ingen lön alls
Tjänsterna för handikappade fås oftast endast med ett läkarintyg (lääkärintodistus).
Rumänska
På FöretagsFinlands telefontjänst får du information, handledning och rådgivning kring start av företagsverksamhet och de offentliga företagstjänsterna.
som har rösträtt i presidentval och
JA: alla leksaker och utrustning som fungerar med el eller batteri
Det lönar sig också att ta med meddelandet om rösträtt.
Om du misstänks för ett brott
Rådgivningen är avgiftsfri.
Socialväsendet bekräftar ett avtal om barnens boende, vårdnad, umgängesrätt och underhållsbidrag.
En utredning över grunden för att den person som ansöker om familjeförening vistas i Finland.
Läkaren diskuterar minnesproblemen med patienten och eventuellt också med dennes närstående och gör ett enkelt minnestest.
Ring inte nödnumret om det inte är fråga om en nödsituation.
Stadsteaternfinska
När beslutet om upplösning har fattats och tillgångarna överlåtits görs en anmälan om upplösning av föreningen till registerstyrelsen.
Skriftlig begäran kan lämnas in till vilken magistrat som helst.
Jämför läkarpriserfinska _ engelska
Edupoli ordnar yrkesutbildning för vuxna.
Hyresboende
Finska för kvinnorfinska
Läs mer om dagvård på InfoFinlands sida Dagvård.
Du hittar kontaktuppgifterna via din hemkommuns webbplats.
Du kan bli intagen på sjukhus med en läkarremiss.
De anställda inom uppsökande ungdomsarbete hjälper med att klara upp den ungas livssituation, hantera praktiska ärenden, såsom besök hos olika myndigheter, och ger personlig handledning enligt den ungas önskemål.
Om du har hemkommun i Finland kan du boka tid för en urologisk undersökning på din egen hälsostation.
De vanligaste hjälpmedlen för synskadadefinska
Vid vårt vetenskaps- och konstuniversitet fås utbildning och idkas forskning inom pedagogik, turism och affärsverksamhet, juridik, konstindustri och samhällsvetenskaper.
Graviditetstest kan köpas till exempel på apoteket.
Du kan få ett tillstånd för högst ett år.
Stadens hyresbostäder
Information för bostadslösafinska _ svenska _ engelska
Utöver modersmålsprovet kan du skriva prov i följande andra ämnen:
Julen
Tillsammans kan ni fundera på vilken sorts stöd som skulle passa just dig.
Om du hittar en arbetsplats, kan du börja arbeta genast.
du är medborgare i EU, Schweiz eller Liechtenstein och du har registrerat din uppehållsrätt i Finland
Därefter flyttas eleven till en vanlig klass.
Även stora mataffärer säljer graviditetstest.
Styrelsens storlek kan föreskrivas i stadgarna.
I den offentliga sektorn (arbetsgivaren är en kommun eller staten) ingås tjänstekollektivavtal eller allmänt kommunalt tjänste- och arbetskollektivavtal.
Hjälp med familjeåterföreningen
Om du behöver ett skattekort eller skattenummer kan du besöka Västra Finlands skattebyrå.
Enligt lag får hyresvärdar inte diskriminera någon till exempel på grund av etniskt ursprung, religion eller medborgarskap när de väljer hyresgäster.
Man kommer punktligt till arbetet på den avtalade tiden.
Alla som bor eller vistas i Finland måste följa Finlands lagar.
Du kan anlita en tolk när som helst om du bokar tolken och betalar kostnaderna själv.
Vid fastställande av skäliga boendekostnader beaktas
I stora städer och deras näromgivning finns en välfungerande lokaltrafik.
Sköta ärenden på Internetfinska _ svenska _ engelska
Om du har en rättsskyddsförsäkring (oikeusturvavakuutus), som ersätter dina utgifter, kan du inte få offentlig rättshjälp.
utfärdar personbeteckningar för personer bosatta i Finland,
InfoFinland-redaktionen sköter uppdateringen av uppgifterna i avsnitten Flytta till Finland, Livet i Finland och Information om Finland samt uppgifterna om Helsingfors, Esbo, Vanda och Grankulla.
Läs mer: Att grunda ett företag.
Du studerar alltså inte vid arbets- och näringsbyrån utan vid den läroanstalt som ordnar kursen.
Ministerierna bereder de ärenden som regeringen fattar beslut om.
I svenskan finns också många lånord från till exempel franskan.
Arabisktalande klienter: 020 634 4902
Hyresvärden kan ange ett konto på vilket du sätter in hyresdepositionen.
Du hittar en lista över kurserna i finska på medborgarinstitutets webbplats.
Observera att samtalspriset ändå alltid beror på vilket land du ringer till.
Läs mer: Kulturer och religioner i Finland.
Utbildning på andra stadiet är oftast kostnadsfri för studeranden.
Du ingår ett elavtal genom att ringa ett elbolag och uppge ditt namn och din nya adress.
Tfn 0800 97899
Grundandet av en förening sker i praktiken i tre steg:
Utvecklingsstörda och arbetefinska
Övriga förmåner för pensionärer
Mottagare av statsförvaltningens språkexamina, finska språketfinska _ svenska
linkkiDroglänken:
Du kan vara pappaledig samtidigt som barnets mor är mamma- eller föräldraledig.
Tfn 045 639 6274
Skatteåterbäring och kvarskatt
pass eller
du har ett gemensamt barn tillsammans med din sambo (då uteblir kravet på gemensamt boende under två års tid)
Stadens ungdomstjänster driver sju ungdomsgårdar runt om i Karleby.
På webbsidorna för Föreningen för mental hälsa i Finland hittar du information om
Du måste också själv ansvara för levnadskostnaderna i Finland.
Betala bolagsvederlag och eventuellt även finansieringsvederlag för bostadsaktiebolagets lån till bostadsaktiebolaget.
barnets far avled innan barnet föddes, barnet föds utom äktenskap i Finland och faderskapet fastställs.
Motionsföreningfinska
Du kan även be om hjälp om du inte vet vilken myndighet du ska kontakta.
Tfn (09) 310 13030
För äldre personer ordnar kommunerna hemvård (kotihoito) som omfattar hjälp med vardagssysslor och sjukvård i hemmet.
Tillståndet är i kraft ett år.
Lag om jämställdhet mellan kvinnor och män
Om du har arbetat i sammanlagt tre år eller mindre, kan du få grunddagpenning i högst 300 dagar.
anpassningsträning
stöd för närståendevård av personer under 65 och arbetsverksamhet.
Om uppgifterna om en utländsk maka eller make inte kan kontrolleras i befolkningsdatasystemet måste personen lämna ett intyg från myndigheterna i sitt eget land för prövning av äktenskapshinder till magistraten.
En förälder till ett barn under 21 år
Om den avlidne har bott eller arbetat utomlands en lång tid innan flytten till Finland, kan de efterlevande även ha rätt till familjepension från det landet.
I staden finns flera cykelleder och vägar som lämpar sig för cykling.
Du kan få rehabilitering till exempel vid en rehabiliteringsinrättning (kuntoutuslaitos).
När du har inreseförbud kan du inte besöka Finland eller något annat Schengenland.
Om äktenskapet har ingåtts utomlands måste man uppvisa ett legaliserat och översatt vigselintyg i magistraten för registrering.
betjänar utomlands bosatta finländare när de behöver sköta ärenden med finska myndigheter, till exempel ansöka om nytt pass
Om du ska vistas i Finland mer än 90 dagar och är EU-medborgare, måste du registrera din uppehållsrätt.
Enligt lagen om likabehandling (Yhdenvertaisuuslaki) får ingen diskrimineras på grund av ålder, etniskt eller nationellt ursprung, nationalitet, språk, religion, övertygelse, åsikt, hälsotillstånd, funktionshinder, sexuell läggning eller av någon annan orsak som gäller hans eller hennes person.
De vanligaste alternativen efter grundskolan är gymnasium och yrkesutbildning.
Ansökan kan göras elektroniskt via stadens webbplats eller med en pappersblankett.
Du kan skriva ett testamente (testamentti), d.v.s. en skriftlig utredning över vem som ska ärva din egendom efter din bortgång.
Den centrala målsättningen är att producera verksamhet som samtidigt är uppfostrande och intressant för de unga, som stöder deras utveckling och uppväxt och som stärker deras samhälleliga delaktighet.
att alltid när det är möjligt bli tillfrågad om sitt medgivande innan behandlingen påbörjas
Hyresbostäder för studerandefinska _ svenska _ engelska
Både ungdomar och vuxna kan studera vid gymnasiet.
Om preventionen misslyckades eller om du glömde att använda preventivmedel kan du köpa ett akut p-piller på apoteket utan recept.
Den unga kan ansluta sig till ett trossamfund eller utträda ur ett trossamfund med föräldrarnas skriftliga tillstånd
Kurser i finska och svenska språketfinska _ svenska _ engelska
Riksdagsval
Kansankatu 8 (vån. 2)
I Finland är kroppsaga på barn (våld i syfte att straffa) förbjuden i lag.
du är gift eller annars i ett nära familjeförhållande till en person som redan bor stadigvarande i Finland.
Service på engelska 0295 020 713
MoniNet, centret för mångkulturell information och verksamhet
Omfattas du av den sociala tryggheten och kan du få bidrag?
Från kunskapscentret får du även rådgivning på telefon eller via e-post när du behöver råd om fostran av barn eller relationerna i familjen.
Hos familjerådgivningen eller vid familjecentret får barn, unga och familjer hjälp med problem som rör fostran av barn och barns utveckling.
När man talar är det oartigt att höja rösten, speciellt på allmänna platser.
Problem med uppehållstillståndet
familjemedlem
Chefen ger den anställda arbetsuppgifter och förväntar sig att den anställda själv fattar beslut om detaljerna i arbetets utförande.
Du hittar information om kurser i finska till exempel hos medborgarinstitut, arbetarinstitut, universitet och sommaruniversitet.
Lapplands TE-byrå
Läs mer:
Ett barn under tre år kan vara i kommunal dagvård på deltid under tiden för flexibel vårdledighet.
Du kan kontakta skyddshemmet även när en familjemedlem har hotat dig med våld.
Om du bor i Finland kan du ha rätt till moderskapsunderstöd (äitiysavustus).
På basis av bedömningen beslutas om boendet är stadigvarande eller inte.
Där hittar man böcker på över 60 olika språk.
Permanent uppehållstillstånd kan eventuellt inte beviljas om:
Beslutsfattande och påverkan
Information om att ansöka om asyl hittar du på InfoFinlands sida Till Finland som asylsökande.
I Rovaniemi finns kommunala daghem och privata daghem.
För att du ska kunna få uppehållstillstånd måste du ha tillräckliga medel för ditt uppehälle.
Hos en privat hyresvärd kan det gå snabbt att få en bostad, men hyran kan vara högre än i stadens hyresbostäder.
Också många företag erbjuder tolktjänster.
kriser
ingen aptit
Om du är en före detta finsk medborgare kan du på denna grund få uppehållstillstånd i Finland.
Tjänsten Miehen Linja (Miehen Linja) är en tjänst som hjälper män, som har utsatt sin partner för våld.
Du behöver inte lämna dricks, men du kan göra det om du vill tacka för en speciellt bra service.
Privat tandvård och ersättningarfinska _ svenska _ engelska
Observera att inloggning till Wilma sker på olika adresser i olika städer.
Brott
Om du är intresserad av adoption, fråga om råd vid socialbyrån i din hemkommun.
Du kan endast söka asyl för dig själv.
Du kan avlägga allmän språkexamen (yleinen kielitutkinto) i finska eller svenska i Esbo.
Knektbrovägen 4
Efter detta bor du i bostaden på hyra och betalar hyra varje månad.
Läs mer på InfoFinlands sida Hemkommun i Finland.
En moder kan bli moderskapsledig redan 31–50 vardagar innan det beräknade förlossningsdatumet.
linkkiNärståendevårdare och Vänner -Förbundet rf:
Kontakta oss om du behöver råd och hjälp i vardagen, vill lära dig finska eller frivilligarbeta, delta i utflykter och evenemang eller utöva fritidsintressen.
Migrationsverket handlägger din ansökan och fattar ett beslut.
Peluuri finns även på internet.
VALMA-utbildningen räcker ett läsår.
Parlamentet har 754 ledamöter och tretton av dem har valts i Finland.
Ansök om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland:
Därtill ordnar Vanda stad filmvisningar.
Elarbeten som du får göra självfinska _ svenska _ engelska
Syftet med serviceplanen är att reda ut vilken handikappservice du behöver.
När du har en bostad är det bra att ta en hemförsäkring.
Migrationsverkets närmaste tjänsteställe finns i Helsingfors:
Arbetstid
På nätet hittar du finskakurser på många olika nivåer.
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lö-sö kl. 8–21.
I Grankulla beslutas ärenden av stadsfullmäktige.
Civil begravningfinska _ svenska _ engelska
Kom ihåg att meddela din arbetsgivare om moderskapsledigheten senast två månader innan den börjar.
Undervisningen sker oftast kvällstid.
Grundläggande utbildning för vuxna invandrarefinska _ engelska
Makarna kan ansöka om skilsmässa tillsammans eller också kan den ena maken göra det ensam.
Läs mer: Mental hälsa.
För att familjemedlemmarna ska kunna få uppehållstillstånd, krävs det i vissa fall att flyktingen har en tillräcklig inkomst för att försörja sina familjemedlemmar i Finland.
Grammatiken Iso suomen kielioppi på nätetfinska
Grundläggande utbildning för invandrarefinska
Du behöver en finländsk personbeteckning och ett finländskt skattekort.
Vilken som helst av vårdnadshavarna kan vara föräldraledig.
Läs mer: Flytta till Rovaniemi
Finlands område var Sveriges buffert österut och gränserna drogs om flera gånger i samband med olika krig.
finns information om familjer som bildas av samkönade par.
Målet med rehabiliteringen är att stöda dig och dina närstående så att du kan föra ett aktivt liv.
Du behöver ha en personbeteckning när du sköter ärenden med myndigheter.
Invandrartjänster
Yrkesinriktad rehabilitering ordnas av arbetspensionsanstalter (työeläkelaitokset) och FPA (Kela).
Migrationsverket ersätter resekostnaderna endast i det fall att familjemedlemmen reser till Finland på en resa som arrangeras av Finlands Röda Kors och Internationella organisationen för migration.
Om du har hemkommun i Helsingfors, kan du använda de offentliga hälsotjänsterna.
Om du saknar pass eller ett identitetskort för utlänningar kan du ta reda på vilken typ av identitetshandling banken kan godta.
linkkiArbets- och näringsbyrån:
linkkiFinlands Näringsliv:
Du kan framföra en begäran om en inledande kartläggning av din situation t.ex. till arbets- och näringsbyrån eller socialbyrån i din kommun.
Du kan också boka tid vid preventivrådgivningen (ehkäisyneuvonta) antingen ensam eller tillsammans med din partner.
I riksdagsval är landet indelat i valkretsar.
En arbetstagare som är medlem i en arbetslöshetskassa betalar en medlemsavgift till arbetslöshetskassan när han eller hon förvärvsarbetar.
Ett samboförhållande är ett förhållande där ett par lever tillsammans utan att vara gifta.
Utländska medborgares bankärendenfinska _ engelska
Handläggning av asylansökan
När brottmålet övergår till domstolen, hålls en rättegång i tingsrätten.
Din sambo som du har bott tillsammans med i minst två år eller med vilken du har gemensam vårdnad om ett barn
En del fritidsaktiviteter är avgiftsbelagda men det finns också tillgång till gratis aktiviteter.
Grunddagpenningen beviljas och utbetalas av Fpa.
Mer information om uppehållstillstånd för arbetstagare och företagare hittar du på sidan Arbeta i Finland och Till Finland som företagare.
Om du avser att bo i Finland längre än tre månader, måste du registrera din uppehållsrätt hos Migrationsverket (Maahanmuuttovirasto).
du har ett uppehållstillstånd som ger dig rätt att arbeta i Finland
I Vanda finns finskspråkiga och svenskspråkiga grundskolor (peruskoulu).
Stäng alltid kranen till tvätt- och diskmaskinen när du inte använder dem.
Att röra sig i naturen är en traditionell och populär form av avkoppling för finländarna under alla årstider.
Evenemangskalenderfinska
Läs mer: Museer.
Mer information om likabehandling hittar du på InfoFinlands sida Jämställdhet och likabehandling.
värnplikt för män (armé eller civiltjänstgöring)
Finansiering av studierna
Nära vänner eller släktingar kan även hälsa på varandra genom att krama om varandra.
I Dickursby finns en ortodox kyrka.
Du kan söka en tolk eller översättare med hjälp av sökfunktionen på Finlands översättar- och tolkförbunds webbplats.
Handikapporganisationer
linkkiBarnombudsmannen:
Du kan även fråga din lärare i finska.
De flesta av FPA:s förmåner är sådana att du har rätt till dem endast om du flyttar ditt stadigvarande boende till Finland eller om din anställning varar i minst fyra månader.
Fortbildning ordnas bland annat av läroanstalter, fackförbund och Institutet för Yrkenas befrämjande.
I Finland ges dagvård, förskoleundervisning och grundläggande utbildning vanligtvis på finska eller svenska.
Information om att leva i ett samboförhållande i Finland hittar du på InfoFinlands sida Samboförhållande.
Rehabilitering som ordnas av FPA
linkkiHelsingfors Företagare:
Mer information får du vid socialbyrån i din hemkommun.
kan du ha rätt till integrationsutbildning som ordnas genom TE-byrån.
Förändringen kan påverka webbplatsens funktionalitet.
På vissa orter kan även socialbyrån (sosiaalitoimisto) eller församlingarna hjälpa.
I tillgången till dagvårdstjänster är målet att uppfylla närserviceprincipen för varje barn.
Du kan också boka tid till läkare på en privat hälsostation.
Om ni har ingått ett avtal om umgänget, men den förälder som bor med barnet inte följer avtalet kan den förälder som bor annanstans kontakta barnatillsyningsmannen i kommunen.
Landhöjningen har varit en central faktor i Karlebys historia.
linkkiFöretagarnas Arbetslöshetskassa i Finland:
Språkkaféerfinska _ engelska _ ryska
rehabilitering för gravt handikappade
Om du tar tillbaka köpeanbudet kan du bli tvungen att betala säljaren böter eller en handpenning.
Läs mer: Förskoleundervisning
Förmånshandläggare
Vid behov kan hälsovårdaren ge remiss till läkare.
Köpa bostad
Man kan också bo tillfälligt i ett familjehem.
Läs mer på InfoFinlands sida Registrering som invånare.
Utkomststöd
Omatila (Omatila) hjälper dig om du har blivit utsatt för närståendevåld eller våld inom familjen.
MoniNet
Patientombudsmannens tjänster är tillgängliga på alla ställen där hälsovårdstjänster tillhandahålls, till exempel på hälsostationer, sjukhus, privata läkarstationer, åldringshem och vårdanstalter för handikappade.
Ungdomarna studerar vid daggymnasiet (päivälukio) eller distansgymnasiet (etälukio), vuxna studerar ofta vid vuxengymnasiet (aikuislukio).
Information om lokala tjänster
Karleby verksamhetsställe
Mer information om tjänsterna för äldre hittar du på Vanda stads webbplats.
Stadens tjänster för arbetssökandefinska _ svenska _ engelska
Om den ena föräldern är hemma, beror rätten till småbarnspedagogik på hemkommunen.
Rådgivning i uppehållstillståndsärenden
Läs mer: Att grunda ett företag i Finland.
Du måste ansöka om ditt första uppehållstillstånd innan du kommer till Finland.
Om du har arbetat i sammanlagt tre år eller mindre, kan du få inkomstrelaterad dagpenning i högst 300 dagar.
Hyresvärden får endast beträda bostaden i vissa undantagsfall, till exempel för att övervaka reparationer i bostaden eller visa bostaden för köpare.
I Esbo finns tre högskolor:
Information om beskattningen av företag och företagarefinska _ svenska _ engelska
Med uppsägningstid avses den tid som avtalet är i kraft efter att det sagts upp.
Det gäller till exempel äktenskapsintyg som utfärdats i USA.
På 1400-talet blev Esbo en självständig socken med många byar.
Får man göra så?
Delta i stämmor och på dem påverka det som händer i bostadsaktiebolaget.
Stadens hyresbostäderfinska _ svenska _ engelska
rådgivning om rehabilitering
Besök till exempel din egen hälsostation för en hälsoundersökning.
Om flera personer har medverkat ska man i sluttexterna ange en ansvarig person som fyllt 15 år.
Tfn: 040 70 46 818
Hur många besökare webbplatsen har
I Finland uppfattas ögonkontakt som uppriktighet och ärlighet gentemot den andra.
Du kan inte söka till ett vuxengymnasium i den gemensamma ansökan.
Lämna till exempel ditt telefonnummer och din adress till TE-byrån och ange hur länge du ämnar vistas på resmålet.
Du kan även fylla i anmälan på magistraten.
Du kan fråga om tolktjänsterna närmare till exempel vid Esbo stads invandrartjänster.
Information om barnskyddslagenfinska _ svenska _ engelska _ ryska _ franska _ somaliska _ persiska _ arabiska _ kurdiska
Tidsenliga intyg
På en stämma kan du rösta om olika saker och kräva att ett ärende tas upp för behandling på stämman.
I Esbo finns flera museer.
Läs mer: Boende.
Du kan också söka ersättning från FPA även i efterhand.
Läs mer: Beskattning
Läs mer: Tandvård.
Återvinningsstationerfinska _ svenska _ engelska
Enligt den överenskomna tidtabellen kommer kärnkraftverket att producera el år 2024.
Kulturer och religioner i Finland
Mottagning /Ullava
Täck inte över dem.
Du kan boka tid vardagar kl. 8–16 på numret 09 816 31300.
linkkiMIELI Psykisk Hälsa Finland rf:
talförståelse
Läkaren bedömer din hörselskada och därefter kan du få hjälpmedel i form av medicinsk rehabilitering.
Du kan få kommunal rehabilitering om du har hemkommun i Finland.
Om du insjuknar akut eller råkar ut för en olycka får du akut sjukvård även om din hemkommun inte är Vanda.
Mete (med metspö) och pimpelfiske omfattas, med vissa undantag, av allemansrätten och du behöver inte skaffa dig ett fisketillstånd för dessa.
Högskolor
TE-byråerna i Östra centrum och Böle gör inledande kartläggningar.
Du kan söka till ett universitet om du har avlagt en finländsk studentexamen, en utländsk examen som motsvarar studentexamen eller en yrkesinriktad slutexamen. Sök till ett universitet i den gemensamma ansökan till högskolor.
Information för nordiska medborgarefinska _ svenska _ engelska _ norska
Utbildnings- och arbetslivsguide för unga(pdf, 26 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska
Filmklipp om motionsalternativfinska _ engelska _ somaliska _ arabiska
Om du har problem i ditt äktenskap eller parförhållande kan du kontakta familjerådgivningen.
När du använder den elektroniska blanketten behöver du finländska nätbankkoder.
Du hittar information om den finländska arbetskulturen på InfoFinlands sida Den finländska arbetskulturen.
Om du har en anställning kan du tala med företagshälsovårdens läkare om sådant som rör den mentala hälsan.
Albertsgatan 25
Antalet intjänade semesterdagar beror på anställningstiden i år och när anställningen har börjat.
Kamrersvägen 3 B
Den ena maken kan inte utan den andra makens tillstånd sälja familjens gemensamma bostad eller tillhörande lös egendom, såsom möbler.
Växel 029 55 39391
Patienternas rättigheter gäller offentliga och privata hälsovårdstjänster samt hälsovårdstjänster till exempel för åldringar och handikappade.
Mer information får du på Utbildningsstyrelsens webbplats.
Mer information om kommunens rehabiliteringstjänster får du vid din egen hälsostation.
Den beräknas oftast på basis av de arbetsinkomster som bekräftats i beskattningen.
Om en ung har problem med alkohol, droger eller spelande, kan hen få hjälp vid ungdomsstationen.
På valet av företagsform inverkar bland annat antalet grundare, behovet av kapital, fördelningen av ansvar och bestämmanderätt, finansieringen och beskattningen.
12 år
Det är möjligt att vårdutgifterna tas ut av dig i efterskott.
Adress: Vasagatan 5
Om högsta förvaltningsdomstolen beviljar besvärstillstånd, behandlar den besvären.
En kvinna behöver inte sin makes eller sina föräldrars tillåtelse för att arbeta eller studera.
När du har bokat tid till tandvård, är det viktigt att komma i tid.
Kom överens om anställningsavtalets innehåll med arbetsgivaren.
Nämnden behandlar ansökningar som berör diskriminering och den kan förbjuda diskrimineringen.
Med vilka apparater och webbläsare sidorna används
Telefontjänsten har öppet måndag till fredag kl. 9.00–16.15.
Stöd betalas för hyra,vederlag och utgifter för skötseln av bostaden.
Du kan vanligtvis ansöka om ett stipendium samtidigt som du ansöker om en studieplats.
du är finsk medborgare och fyller 18 år senast på valdagen,
Arbetslagstiftningen och kollektivavtalen föreskriver vilka rättigheter och skyldigheter arbetstagare har.
Vårdledigheten kan vara högst fyra dagar.
Om du misstänker att ditt barn eller din ungdom behöver barnskyddets (lastensuojelu) hjälp, ska du kontakta en socialarbetare.
Missbruksproblem hos ungdomar
Läs mer på InfoFinlands sida Bibliotek.
Mer information om legalisering av handlingar får du hos magistraten eller hos ditt lands beskickning i Finland.
tfn 016 3223 412
Du kan söka handikappbidrag hos FPA.
Vissa små elarbeten får du utföra själv, om du kan.
Du kan kontakta rådgivningen om du tror att du har blivit utsatt för diskriminering.
Om du omfattas av den sociala tryggheten i Finland ersätter FPA en del av kostnaderna.
Böcker och annat studiematerial måste man dock köpa själv.
Det riksomfattande servicenumret är 0295 025 500 på finska, 0295 025 510 på svenska, 0295 020 713 på engelska och 0295 020 715 på ryska.
Statskontorets tjänsten Medborgarrådgivning hjälper medborgarna att snabbt och smidigt hitta rätt myndighet eller elektronisk myndighetstjänst.
Om du får ett jobb kan du börja arbeta direkt.
Din makes/makas inkomster inverkar inte på din skatteprocent.
Ett tidsbundet avtal kan hävas endast av mycket vägande skäl.
Du kan söka dessa företag till exempel med sökmotorer på Internet.
Den partiella sjukdagpenningen (osasairauspäiväraha) är avsedd för 16–67-åriga heltidsarbetande anställda eller företagare som omfattas av den sociala tryggheten i Finland.
Söka asyl
Vid Österbottens TE-byrå (arbets- och näringsbyrå) får du hjälp med att hitta en arbetsplats.
Till exempel ska en badrumsrenovering alltid meddelas i förväg.
Den finska personbeteckningen är en nummerserie med elva siffror som bildas baserat på ditt födelsedatum och ditt kön.
Fiske och jaktfinska _ svenska _ engelska
Invandrartjänsterfinska _ svenska _ engelska
Varken du eller din sambo får vara gift med någon annan.
Dessutom ska minst två vittnen som har fyllt 15 år vara på plats.
Esbo tillhör samkommunen Helsingforsregionens trafik HRT (HSL), som ordnar kollektivtrafiken i huvudstadsregionen.
Trots att du inte har uppehållstillstånd kan du börja arbeta när du vistats i sex månader i landet.
Anmälan till skolanfinska _ svenska _ engelska
Stödcentret Hilma för handikappade invandrare
Läs mer: Föreningar.
Om du inte har hemkommun i Finland och inte heller någon annan grund ger dig rätt att utnyttja de offentliga hälsovårdstjänsterna i Finland måste du betala ett pris som motsvarar de faktiska kostnaderna för dessa hälsovårdstjänster.
Ett rasistiskt brott kan vara till exempel våld, ärekränkning, diskriminering, hot, trakasserier eller skadegörelse.
Rådgivningen hjälper dig att fylla i ansökan.
Du kan också söka hjälp för en familjemedlem eller en vän.
Det lönar sig att söka hjälp, om du har något av följande symptom:
Kurserna är avgiftsbelagda.
Kopian kan pålitligt vidimeras av den myndighet som utfärdat handlingen eller notarius publicus i det land där handlingen utfärdades.
Nylands TE-byrå (TE-toimisto) erbjuder mångsidiga tjänster för personer som funderar på att starta eget och dem som är på väg att starta eget.
Televisionen i Finlandengelska
Du kan fråga mer om tjänsterna vid enheten för socialarbete i ditt bostadsområde.
På InfoFinlands sida Familjer med en förälder finns information om hurdant understöd den vårdnadshavare som bor med sitt barn kan få om föräldrarna inte bor tillsammans.
Hyreshandboken(pdf, 1,11 MB)finska _ svenska _ ryska _ franska _ somaliska _ arabiska
+358 (0)29 497 151 (svenska)
är 17–64 år gammal
Utlåtanden om utländska yrkesexamenfinska _ svenska _ engelska
Läs mer om fortsatta studier på InfoFinlands sidor Universitet och Yrkeshögskolor.
Socialservicecentret
Du kan avlägga studier vid öppna högskolan fastän du får arbetslöshetsersättning (työttömyyskorvaus).
Du behöver inte uppge ditt namn då du ringer.
– Du kan även lyfta fram dina intressen.
Om du behöver stöd eller är orolig för barnet är det bäst att i god tid be om råd till exempel vid den egna kommunens socialtjänst.
Mellersta Österbottens utbildningskoncernfinska _ engelska
Undersökning av bröstcancer görs på kvinnor i åldern 50–69 år ungefär vartannat år.
Läs mer: Barn vid skilsmässa.
För vissa arbetsuppgifter behöver du inte ett uppehållstillstånd för arbetstagare, men du behöver dock ett uppehållstillstånd som beviljas för vissa uppdrag.
Arbetslöshetsersättning
Valet förrättas vart femte år.
När du söker en studieplats krävs inte nödvändigtvis erkännande av examen.
engelska 029 497 050
Du kan bli tvungen att vänta länge på en bostad.
Till den finländska julen hör många slags festmat, såsom julskinka, rosoll som är en rödbetssallad, olika slags lådor, julstjärnor och pepparkakor.
Uppehållstillstånd för arbetssökande kan beviljas för högst ett år.
TE-byrån betjänar på internet via sidan E-tjänster (Oma asiointi).
Behovet av närståendevård för personer under 65 år bedöms inom handikapprådgivningen.
Färdighetsnivåerna i allmänna språkexaminafinska _ svenska _ engelska
Om din inkomst har ökat kan du söka sjukdagpenning på basis av arbetsinkomsten under de senaste sex månaderna.
I den grundläggande utbildningen ges alla vitsord av läraren.
Kontakta mödrarådgivningen direkt i början av graviditeten.
Du får blanketten från magistraten eller på magistratens webbplats.
linkkiRegnbågsfamiljer:
Rörelsehandikappade
Kom med och bygg framtidens InfoFinland!
Försäkringens självrisk får inte överstiga 300 euro.
Barnrådgivningens arbete omfattar barn under skolåldern och deras familjer.
Ansök om studieplats
I annat fall förfaller ärendet.
Om denna stat inte tillåter flerfaldigt medborgarskap kan du förlora ditt nuvarande medborgarskap när du får finskt medborgarskap.
Mer information hittar du på Migrationsverkets webbplats.
uppehållskort;
Föreningar
Om du är under 30 år kan du få informations-, rådgivnings- och handledningstjänster på Rovaniemi stads navigator.
ett kombinerat efternamn som har bildats av föräldrarnas efternamn.
Daghem och skolor gör sitt för att ordna motion men detta är inte deras huvudsakliga uppgift.
Om du misstänker att du har blivit utsatt för diskriminering, kan du kontakta Brottsofferjourens rådgivning för att motarbeta diskriminering.
Grunden för din vistelse kan ändras till exempel om du får en arbetsplats i Finland eller gifter dig med en finsk medborgare eller en person som har kontinuerligt eller fortsatt tillstånd i Finland.
År 2002 införde Finland bland de första EU-länderna EU:s gemensamma valuta, euro, och gav därmed upp sin egen valuta.
Norrsken
bostadsort
FPA kan delvis ersätta resorna till rehabiliteringen.
Ett lätt sätt att komma igång är till exempel genom att delta i skolans eller läroanstaltens elevverksamhet.
Erkännande av examen är avgiftsbelagt och söks hos Utbildningsstyrelsen.
Om du insjuknar måste du själv betala läkar- och sjukhuskostnaderna.
Olika regioner i Finland har olika matkulturer.
Information om kyrklig vigselfinska _ svenska _ engelska
I Finland börjar den grundläggande utbildningen det år då barnet fyller sju år.
Om du är studerande kan du ansöka om en hyresbostad via Helsingforsregionens studentbostadsstiftelse HOAS (Helsingin seudun Opiskelija-asuntosäätiö HOAS).
På InfoFinlands sida Ring och fråga om råd hittar du mer rådgivningstjänster.
tillfälligt vistas på marker där det är tillåtet att röra sig enligt ovan. Du kan till exempel tälta relativt fritt bara du håller ett tillräckligt avstånd till andras bostäder.
Att följa ordningsreglerna i ditt bostadsaktiebolag om du bor i ett höghus eller ett radhus.
Läs mer: Dödsfall.
Hjälp med penningspelproblemfinska
Diskrimineringsombudsmannen är en myndighet vars uppgift är att främja likabehandling och ingripa i diskriminering.
Äldre människor
Utöver den finns det flera kommersiella tv-kanaler i Finland, till exempel MTV3 och Nelonen.
linkkiFörbundet för mödra- och skyddshem:
På så sätt säkerställer du att du inte ställs ansvarig för fel som du inte har orsakat.
Fråga mer om detta vid beskickningen för ditt eget land.
Du kan få studielån också när du fortbildar dig (täydennyskoulutus) som vuxen.
Det finns en biograf i Grankulla.
Läs mer: Trafiken.
I Vanda finns många privata läkarstationer som även tar hand om barn.
Adress: Hermanstads Strandväg 12 A, vån. 4
Det kan exempelvis vara avgångsbetyg från finsk grundskola.
Du får information om hur du köper en bostad på InfoFinlands sida Köpa bostad.
Ryssland gjorde området som erövrats till Finlands autonoma storfurstendöme.
Du kan gå till en privat tandläkare även om du inte har rätt att använda den offentliga hälsovårdens tjänster.
Esbos areal är cirka 528 km2, varav cirka 216 km2 är vatten.
FPA:s ersättning kan ibland dras av direkt på det belopp som du betalar vid kassan.
Ett barn kan samtidigt ha både finskt medborgarskap och medborgarskap i ett annat land, om det andra landet godkänner flerfaldigt medborgarskap.
Du hittar kontaktuppgifterna till daghemmen på stadens webbplats.
Det är bra att en gång per år städa bort damm från frysens och kylskåpets bakgaller till exempel med dammsugaren, om möjligt.
De tre månaderna räknas från den dag då din maka/make/sambo/partner delgivits beslutet.
Finland lyckades dock skapa goda relationer till Sovjetunionen, bibehålla sitt demokratiska system och öka handeln också med västländerna.
Till exempel ligger Helsingfors-Vanda flygplats i Vanda.
Om du flyttar till Finland för att studera kan du inte få studiestöd.
I de flesta situationerna bedömer arbetsgivaren, läroanstalten eller högskolan vilken behörighet och kompetens din utländska examen ger.
den ena föräldern eller båda föräldrarna har hemkommun i Finland eller
Flera kultur- och motionslokaler möjliggör varierande former av hobbyverksamhet.
företagsfinansiering
Läs mer: Högskoleutbildning.
Make eller maka till en finsk medborgarefinska _ svenska _ engelska
Lapplands TE-byrå betjänar kunderna per telefon måndagar, onsdagar, och torsdagar kl. 8–16.15 samt tisdagar och fredagar kl. 9–16.15 på numret 0295 039 501
Beskickningen kan bevilja dig ett nytt pass om ditt pass har gått förlorat eller stulits.
Problem med den mentala hälsan
Ditt permanenta eller tidsbegränsade uppehållstillstånd återkallas om
Trafikförsäkringen tecknar du hos ett försäkringsbolag.
Olika konstarter är musik, bildkonst, dans, teater och cirkus.
Lapplands skogsmuseumfinska _ engelska
Avgiften gäller lägre och högre högskolestudier på engelska.
Akutmottagningen vid Lapplands centralsjukhus
linkkiInternationella föreningen i Håkansböle:
För att du ska kunna söka en hyresbostad hos staden, ska du ha uppehållstillstånd för minst ett år.
Det finns även andra stödformer för nya företagare.
På InfoFinlands sida Problematiska situationer i Esbo hittar du uppgifter om vart du kan vända dig i Esbo för att få hjälp vid barns och ungas problem och problem i familjen.
och om du på grund av din skada behöver hjälp av en tolk
Information om undervisning i elevens eget modersmål och religion får du av koordinatoren för undervisningen för olika språk- och kulturgrupper:
Flexibel eller partiell vårdpenning betalas inte för vård av ett barn som fyllt tre, men som ännu inte går i skolan.
När du har hittat en lämplig bostad bör du snabbt bestämma dig om du vill ha den.
Om arbetsgivaren inte ger en redogörelse för de centrala villkoren i arbetet till den anställda kan han eller hon dömas till böter.
Jag har ett tills vidare gällande hyresavtal.
På biblioteket kan du också använda dator.
Om det är snö och is på marken är det också halt.
Tidningen med den största upplagan är Helsingin Sanomat.
Privat läkarstationfinska _ svenska _ engelska
Migrationsverket beslutar om du ska beviljas uppehållstillstånd eller inte.
Samboförhållande, äktenskap och separation
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Om du inte har rätt att använda de offentliga hälsovårdstjänsterna kan du kontakta en privat läkarcentral.
Att studera i Finland
linkkiEvira:
Mer information om studerandehälsovården får du på Studenternas hälsovårdsstiftelses (SHVS) (YTHS) och social- och hälsovårdsministeriets (Sosiaali- ja terveysministeriö) webbplatser.
Skolornas kontaktuppgifterfinska
Om du är av finländsk härkomst eller har en nära kontakt med Finland kan du beviljas uppehållstillstånd i Finland på grund av detta.
För tillnyktrings- och avgiftningsvård debiteras en patientavgift liksom även för korttidsrehabilitering, öppen rehabilitering är gratis.
Tfn 050 571 5860
Hjälp med att dela egendomen
Visa att du har bekantat dig med arbetsgivarens organisation och arbetsuppgiften i förväg och att du har ett äkta intresse för jobbet.
Du kan få startpeng om
Man måste betala skatt för privatvårdsstödet.
Med infödd finsk medborgare avses en person som har fått finskt medborgarskap vid födseln.
Om du är medborgare i något annat land behöver du ett uppehållstillstånd för arbetstagare.
Luckan Integration är en rådgivningstjänst som erbjuder invandrare personlig rådgivning, och ordnar bland annat möten och grupper i anslutning till arbetssökande.
Information om Humanistiska yrkeshögskolanfinska _ engelska
För skattepengarna betalar staten och kommunerna till exempel:
Våld är alltid ett brott i Finland.
Det gemensamma telefonnumret till servicepunkterna är (09) 816 57070 och e-postadressen är info(at)espoo.fi.
Då beställer myndigheten tolken och betalar för tolkningen.
Handläggningen av ansökan är avgiftsbelagd.
I Vanda finns många motionsslingor och naturstigar.
matrester
fiska eller jaga utan de tillstånd som krävs.
Man kan inte lösa in bostaden, men man kan sälja bostadsrätten eller byta till en annan bostad.
Skolhälsovårdaren har hand om skolelevers hälsa.
Tfn 029 553 9391
02701 Grankulla
Parterna döms till skilsmässa även om den andra parten motsätter sig det.
Om du har avlagt högskolestudier utomlands och vill fortsätta dina studier i Finland kan du få information och handledning vid högskolornas tjänster för studerande och SIMHE-tjänsterna.
Jourhjälpen (Päivystysapu) betjänar dygnet runt.
Du får information om dem vid seniorrådgivningen.
Rättigheterna och skyldigheterna enligt Finlands grundlag gäller alla barn som bor i Finland.
Om det behövs ytterligare utredningar för din ansökan kommer detta att meddelas via ditt konto.
Lån
Privat tandvård
I Finland reglerar lagstiftningen den grundläggande utbildningen.
Ta med dig ett officiellt identitetsbevis när du använder hälsovårdstjänsterna.
Till exempel bedömer arbetsgivare i privatsektorn oftast själv huruvida en utländsk examen ger tillräckliga kvalifikationer för uppgiften.
Gymnasieförberedande utbildning för invandrarefinska _ engelska
Sjukhusgatan 3
Vandainfofinska _ svenska _ engelska
Mer information om hjälp för barn i problematiska situationer får du på InfoFinlands sida Var hittar jag hjälp när barn eller unga har problem?
I Finland finns sju Unescos världsarv.
Telefon: 09 310 11111, mån.–tors. kl. 9–16, fre. kl. 10–15
Du kan köpa biljetter på Matkahuoltos verksamhetsställen och webbplats.
linkkiBrahestadsregionens företagstjänster:
Sjukdagpenningens belopp beror på inkomsterna.
Med äktenskapsförord kan makarna utesluta giftorätten i den andras egendom antingen helt eller delvis om de skiljer sig eller om den ena av makarna dör.
Ett bibliotekskort får du gratis på biblioteket.
Stöd för föräldrarfinska
Mer information om arbete och företagande i Finland hittar du på InfoFinlands sida Arbete och entreprenörskap.
Munhälsafinska _ svenska
Ellfolkgatan 5, 68300, Kelviå
Naturen är mycket viktig för finländarna.
En del läkare inom den offentliga hälsovården gör gynekologiska undersökningar.
Alla har skyldighet att vittna inför domstol om de blir kallade.
Varför bostadsrättsbostad?
Om du inte har rätt att använda de offentliga hälso- och sjukvårdstjänsterna, kan du boka tid på en privat läkarstation.
Försäkring för studerandefinska _ svenska _ engelska
Inträdet kostar i snitt fem euro för vuxna och två euro för barn.
Mer information om uppehållstillstånd för företagare hittar du på InfoFinlands sida Bli företagare i Finland.
Stadsfullmäktige är det högsta beslutsorganet i staden.
Dagarna innehåller mycket lek och utevistelser.
Äktenskapsförord kan upprättas före äktenskapet eller under det.
linkkiSopu-arbetet:
Om du behöver brådskande tandvård, ska du ringa tidsbokningen så fort den öppnar kl. 7.30.
På K.H.Renlunds museums webbplats finns mer information om museets tjänster, utställningar samt aktuell verksamhet.
Beslut om utbetalning av förhöjningsdelen fattas av den som betalar arbetslöshetsförmånen, alltså arbetslöshetskassan eller FPA.
Du kan få inkomstrelaterad dagpenning från företagarnas arbetslöshetskassa om du har bedrivit företagsverksamhet och varit medlem i kassan tillräckligt länge innan du blev arbetslös.
På Infobankens sidor hittar du mycket information om tjänsterna på olika orter.
Svenskspråkiga arbetarinstitutet Arbisfinska _ svenska _ engelska _ ryska
Du hittar byrån för ungdomstjänster vid Salutorget, på övervåningen i Monde ungdomsgård.
Förflyttningstillstånd beviljas av besiktningskontor och vissa av Tullens verksamhetsställen.
Vad kan jag göra?
Friluftskartor på Internetfinska _ svenska _ engelska
Du kan anmäla ditt barn till skolan via Internet eller genom att besöka skolan på anmälningsdagen.
Du kan söka bostad samtidigt på många olika områden.
Lokal information
Med stadigvarande boende i Finland avses att du har ditt egentliga hem i Finland och huvudsakligen också vistas i landet.
EES-länderna är Europeiska unionens medlemsländer samt Norge, Island och Liechtenstein.
Offentlig tandvård är gratis för barn under 18 år.
På våren och hösten ligger temperaturerna här emellan.
Anmälan till grundskolan sker vid den skola som anges i ett brev som varje ny elev får hem eller per telefon till skolan.
Föräldrarna anmäler sitt barn till skolan.
Patientföreningar
Familjer som bor i Grankulla kan också söka dagvårdsplats till sitt barn i Esbo, Helsingfors eller Vanda.
Beslutet om att använda tolk fattas av föräldrarna.
Om du är i ålderspension påverkar din arbetsinkomst inte pensionens storlek.
Om du har en finländsk personbeteckning kan du söka hyresbostad hos Helsingfors stad via internettjänsten stadinasunnot.fi.
Fråga mer om omskärelse på rådgivningen, av läkaren på hälsostationen, skolhälsovårdaren eller skolläkaren.
Deltagande i elev- och föreningsverksamhet är ett bra sätt att bidra till att också de unga får sin röst hör då det fattas beslut om sådant som påverkar deras livsmiljö.
Du behöver inte uppge ditt namn när du ringer.
Ansökan kan även skickas till tingsrättens kansli per post eller via e-post.
Bostaden kan vara:
De flesta studerande som bedriver fortsatta studier avlägger doktorsexamen.
Utbildning som rör arbetet
sambo
Översättningsanvisning:
På boendekostnaderna inverkar
Miestentie 3
Kronoby folkhögskolafinska _ svenska _ engelska
Du behöver ett utlåtande från Business Finland som bifaller verksamheten som tillväxtföretagare.
Ett handikappat barn kan få specialundervisning om barnets handikapp försvårar inlärningen.
Allemansrätten
Karleby stadsbibliotek finns i stadens centrum.
Grundläggande rättigheter
Gymnasiestudierna är mer teoretiskt inriktade än yrkesutbildning.
Du har bott i Finland tillräckligt länge.
Riksdagen (eduskunta) stiftar lagarna i Finland och beslutar om statens budget.
Lediga tjänsterfinska
Mammorna firas till exempel med presenter och blommor.
om ni har bott tillsammans minst fem år eller
Om du behöver boka en tid till TE-byrån ska du kontakta TE-byrån direkt per telefon eller boka en tid på plats.
Internationellt skydd kan beviljas om personen känner välgrundad fruktan för förföljelse (på grund av ras, religion, tillhörighet till en viss samhällsgrupp eller politisk samhörighet) eller om personen annars är utsatt för verklig fara i sitt hemland eller sitt permanenta bosättningsland.
Du kan ansöka till den grundläggande utbildningens tilläggsundervisning, det vill säga till en tionde klass (kymppiluokka), om du fick grundskolans avgångsbetyg samma år eller året innan, men inte har fått en studieplats på andra stadiet.
Om barnet är i skolåldern kan du kontakta skolpsykologen eller skolläkaren.
Som flyttsaker betraktas till exempel:
Om du flyttar från Finland utbetalas arbetspension från Finland då du går i pension.
Om du vill söka en av stadens hyresbostäder ska du fylla i en ansökningsblankett för hyresbostäder.
Du kan även besöka servicestället In To Finland i Kampen i Helsingfors.
Med en allmän språkexamen kan du påvisa dina kunskaper i finska eller svenska.
Utöver modersmålsprovet måste du skriva prov i minst tre andra ämnen.
Kontaktuppgifter till polisstationernafinska _ svenska _ engelska
Du kan ansöka om utkomststöd hos FPA.
Om du har fått din personbeteckning någon annanstans än vid magistraten och vill ha en hemkommun, måste du även besöka magistraten.
Försök att komma överens om att få mer tid på dig att betala.
Under de tysta timmarna får man inte vara högljudd, till exempel spela på instrument eller lyssna på musik på hög volym, men normalt liv är tillåtet.
En brandvarnare räcker till 60 kvadratmeter.
Webbtjänsten InfoFinland hette tidigare Infobanken.
Enligt Finlands lag har män och kvinnor samma rättigheter.
Läs mer: Diskriminering och rasism.
Fritidsverksamhet för barn och unga
Arbetskraftsutbildning (työvoimakoulutus)
En förening kan till exempel vara ett idrottssällskap, en kulturförening, en vänskapsförening eller en religiös förening.
En del av företagets finansiering kan bestå av en gåva eller ett lån.
Kan jag säga upp den senare?
I Finland ordnar kommunerna tjänster för äldre för att underlätta deras vardag och för att de ska kunna bo hemma så länge som möjligt.
Åren 2017–2020 var statens finansiärer arbets- och näringsministeriet, undervisnings- och kulturministeriet, miljöministeriet, FPA och Skatteförvaltningen.
Hur beräknas skatteprocenten?finska _ svenska _ engelska
I Finland lider 20 % av befolkningen av depression i något skede av livet.
Se till att du har en släckningsfilt hemma.
Du kan inte skicka din ansökning via e-post eller fax.
Om videoklippet/verket innehåller material, vars upphovsrätt innehas av en tredje part, ska upphovsmannen säkerställa att han eller hon har vederbörliga tillstånd till att använda materialet.
Internet
Du kan få arbetslöshetsförmån under studierna, om
Val av tävlingens vinnare och pris
Du kan be om hjälp med att beräkna underhållsbehovet hos barnatillsyningsmannen (lastenvalvoja) i din hemkommun.
När det finns ett avgörande om att ditt boende i Finland är stadigvarande, anses du bo stadigvarande i Finland så länge som
Gymnasium.
är arbetsförmögen och tillgänglig på arbetsmarknaden
Ta också reda på om försäkringar täcker de risker som förknippas med verksamheten.
Ekonomisk rådgivning för företagarefinska _ svenska
Ring nödnumret 112 om det är fråga om en brådskande nödsituation.
Du kan använda samma skattekort hos alla arbetsgivarna.
Prata först med din chef.
Som gäst i ett finländskt hem
Du kan också till exempel kontakta grannmedlingscentret Naapuruussovittelun keskus.
följa lagar och avtal
I Helsingfors finns det lekparker och familjehus, där det ordnas verksamhet för barn och föräldrar som sköter barnen hemma.
linkkiEsbo stad:
Grankulla har cirka 9 600 invånare, varav 60 procent har finska, 36 procent svenska och 4 procent ett annat språk som modersmål.
Webbsidorfinska _ svenska _ engelska _ ryska _ kinesiska
En del företag som tillhandahåller flyttservice sköter också flytt från ett land till ett annat.
När du kommer till jourmottagningen ska du ta en kölapp, såvida du inte har en bokad tid.
Hälsovård för papperslösa
En invandrare som har bott tillräckligt länge i Finland kan få pension på grund av sin ålder eller arbetsoförmögenhet.
Telefon: 0295 018 450
I integrationsutbildningen studerar man finska, kommunikationsfärdigheter och mycket annat. För den som flyttar till
Också alkoholdrycker är dyra på restaurang.
I Finland är arbetsgivare skyldiga att ordna förebyggande företagshälsovård för sina anställda.
Kursansökan kan lämnas in via Internet.
Parterna som ingår arbetsavtalet
Läs mer om hjälpmedel och förändringsarbeten på InfoFinlands sida Tjänster för handikappade.
Som heltidsstudier räknas följande:
Hjälptelefoner
Läs mer: Sexuell hälsa och prevention.
I de flesta städer finns en biograf.
Utbytesstudenter kan få studieplats till exempel via Erasmus, Nordplus, FIRST och Fulbright.
Om du har bott eller arbetat i andra EU-länder än Finland eller i något land med vilket Finland har ett socialskyddsavtal, kan du ha rätt till pension från dessa länder.
Vid Esbo stads servicepunkter (asiointipiste) får du mer information om stadens tjänster.
Språket som talas vid träffarna är engelska.
Ibland kan konflikterna mellan olika kulturer skapa problem mellan barnen och föräldrarna.
Längden på skoldagarna varierar i olika årskurser.
Fastighetsskötseln kan göra små reparationer, till exempel reparera en kran eller öppna upp ett avlopp.
Äldre i Helsingfors och deras anhöriga kan kontakta Seniorinfo.
I Helsingfors finns många studiemöjligheter som är öppna för alla.
Folkhögskolor
På denna grund kan uppehållstillstånd beviljas till exempel för en förälder till en myndig (18 år gammal) person.
Du studerar vid en yrkesläroanstalt eller avlägger yrkesinriktade tilläggsstudier
Bil och körning i Finlandengelska
Du kan också boka tid hos en psykiater eller en psykolog vid en privat läkarstation.
Läs mer om finskt medborgarskap på InfoFinlands sida Finskt medborgarskap.
Myndigheten bokar tolken och då får du tolkningstjänsten gratis.
linkkiCentralorganisationen för högutbildade i Finland Akava:
Om föräldrarna inte kan enas om underhållsbidraget kan de få hjälp i form av medling i familjefrågor.
Ungdomsgårdarna är ungdomarnas egna lokaler där de tillsammans med ungdomsledarna kan syssla med sådant som är viktigt för dem.
studierna leder till yrke eller examen
Föräldrapenningperioden varar i cirka sex månader.
Rådgivning för personer som säljer sexuella tjänsterfinska _ engelska
tfn 020 435 4810 Öppet mån–fre kl. 9–16
Studerandes rätt att arbetafinska _ svenska _ engelska
Läs mer på InfoFinlands sida Trafiken i Finland.
Alla klienter inom hälsovården har rätt till likabehandling utan diskriminering.
Du kan söka information om teatrarnas repertoar och tillgängligheten av biljetter och biljettpriserna till exempel på biljettjänstens eller teatrarnas webbplatser.
Asylsamtal
Barnskyddsanmälanfinska _ engelska
Med hjälp av uppföljningen vet vi till exempel följande:
För att kunna ansöka om en hyresbostad hos staden, måste du ha uppehållstillstånd för minst ett år.
linkkiArbets- och näringsministeriet:
linkkiEsbo Företagare:
naturvetenskaper
Om huset värms upp med olja ska du komma ihåg att kontrollera oljemängden.
FPA sköter även de sjukvårdsersättningar som betalas för privat sjukvård.
I Finland har alla företagare bokföringsskyldighet.
InfoFinlands samarbetsavtal
du har vistats utomlands utan avbrott i två år
Välj något annat språk.
Kurser i finska språket vid öppna universitetet
Kontaktuppgifter till servicestället International House Helsinki:
Om du inte har rätt att använda de offentliga hälsovårdstjänsterna, har du rätt att behandlas jämlikt inom den privata hälsovården.
Napapiirin Residuum
För finskt medborgarskap behöver du ett intyg för åtminstone nöjaktiga språkkunskaper.
Också Helsingfors universitets öppna universitet (avoin yliopisto) har verksamhetsställen i Vanda. Där ges undervisning på högskolenivå och fortbildning.
Registrering som invånare.
Innan du ansöker om finskt medborgarskap är det bra att ta reda på om flerfaldigt medborgarskap också är tillåtet i det land där du är medborgare.
På rådgivningsbyrån följs barnets hälsa, tillväxt och utveckling upp och där ges även vaccinationerna.
Man kan komma överens om en prövotid i anställningens början.
Detta förutsätter att du lämnar in en ansökan i ärendet inom ett år efter din flytt utomlands.
Sopsortering och avfallsåtervinningfinska
Information om den förberedande utbildningen får du vid rådgivningen och kundtjänsten vid sektorn för fostran och utbildning eller vid Stadin ammattiopisto.
Om du har ett tills vidare gällande hyresavtal är uppsägningstiden vanligtvis en kalendermånad.
senaste löneintyg
Mer information om öarna och vattentrafiken får du på Helsingfors stads webbplats.
Röda Korset har ett skyddshus för 12–19-åriga unga.
Barn har även rätt att uttrycka sina egna åsikter.
Om du är kund vid arbets- och näringsbyrån kan du också studera svenska som arbetskraftsutbildning.
Den inledande kartläggningen och integrationsplanen kan utarbetas tillsammans med dig antingen på Lapplands TE-byrå eller inom Rovaniemi stads socialservice, till exempel inom de integrationsrelaterade socialtjänsterna
Tjänsten ger dig råd om olika kollektivtrafikförbindelser från ett ställe till ett annat.
När du är gravid:
Om du till exempel oväntat får arbete eller en studieplats kan du ansöka om vårdplats senare.
Registerbeskrivning
Studiepsykologer och skolkuratorer hjälper eleverna i problemsituationer.
I din ansökning ska du motivera varför ditt uppehållstillstånd inte bör återkallas.
Jourmottagningen för barn och unga finns ofta i en separat enhet.
Du kan få studiestöd om
Mer information om Rovaniemi stads idrottstjänster och hälsomotionskalendern hittar du under följande länk:
Besöksförbud
Du kan kontakta den närmaste hälsovårdscentralen (terveysasema), om du har problem med alkohol eller droger.
Läs mer om att grunda ett företag på InfoFinlands sida Att grunda ett företag i Finland.
Unga i åldern 12–19 år kan kontakta Röda Korsets De ungas skyddshus (Nuorten turvatalo).
H-klinikka
– Om du vill kan du även lista dina publikationer eller arbetsprov.
Underhållsförmågan beräknas genom att dra av skatter och övriga obligatoriska utgifter av inkomsterna.
Arbetsgivaren är skyldig att betala lön för sjukledigheten.
Färdtjänst och följeslagartjänstfinska _ svenska
Nedan följer några exempel på yrkesinriktad arbetskraftsutbildning:
Mer information om att ansöka om fortsatt uppehållstillstånd hittar du på InfoFinlands sida Fortsatt uppehållstillstånd.
Via Rovanapa Oy kan du ansöka om en bostad vid Kunta-asunnot Oy.
Det är bra att boka en tid hos beskickningen eller tjänstestället i förväg.
I staden finns också många idrottsmöjligheter.
Diskrimineringslagen definierar vad som är diskriminering.
Om du ärver egendom av en avliden person måste du betala arvsskatt (perintövero) för egendomen.
Webbplatsen asuminen.fifinska _ svenska _ engelska
Om du till exempel flyttar från höghus till egnahemshus behöver du förmodligen en annorlunda försäkring.
högskoleexamen gymnasiestudier eller
Könssjukdomar
För finländarna var det ändå viktigast att ha kunnat bevara landets självständighet.
Grunddagpenning
Trafik
På InfoFinlands sida Bostadsbidrag finns mer information om FPA:s allmänna bostadsbidrag.
Mer information om läkemedel får du på InfoFinlands sida under rubriken Läkemedel.
De flesta finländarna bor i en ägarbostad, alltså i en bostad som de själva äger.
Om du och din sambo är bosatta i olika stater anses gemensamt boende till exempel under semesterresor inte som en tillräcklig grund för beviljande av uppehållstillstånd.
Barnet kan även få undervisning i den egna religionen eller i livsåskådningskunskap i förskolan.
Om du vårdar ditt barn i hemmet och behöver tillfälligt en vårdplats för barnet, till exempel när du ska sköta ärenden, kan du kontakta barnpassningsservicen (hoitoapupalvelu).
Innan äktenskapet ingås ska du skriftligen be om prövning av äktenskapshinder.
Mer information får du på Utbildningsstyrelsens webbplats.
Om du har anlänt till Finland för en kort tid sedan och har barn under skolåldern ska du ta kontakt med områdeskoordinatorn för ditt bostadsområde (aluekoordinaattori).
Små barn behöver inte nödvändigtvis ledd motion, utan det räcker med vanlig lekverksamhet och utevistelser i olika miljöer.
Äktenskapsförordet görs skriftligt. Det dateras och undertecknas.
När du ska fatta beslut om abort får du stöd till exempel av en hälsovårdare eller en läkare vid hälsostationen.
Köpcentret Rinteenkulma
Om din make eller maka bor stadigvarande i Finland, kan du få uppehållstillstånd i Finland på grund av äktenskapet.
Påbyggnadsexamina vid universitetfinska
stället där arbetet utförs
Att bo i en bostadsrättsbostad är ett alternativ till att köpa eller hyra sin bostad.
I vilket land användarna befinner sig
Du kan boka tiden via telefontjänsten eller på FPA:s webbplats.
Om det förekommer våld eller missbruk i familjen ingriper barnskyddets socialarbetare i situationen.
Flyktingsrådgivningen bistår asylsökande juridiskt i asylprocessen.
Du kan även studera flera andra språk, såsom engelska eller franska.
Du ska meddela FPA och arbetspensionsanstalten om du börjar arbeta.
Då kan du välja läkaren själv.
Vi erbjuder allt textinnehåll i InfoFinland via ett öppet programmeringsgränssnitt (API).
Om du är medborgare i ett EU-land, ett EES-land, Schweiz eller i något av de nordiska länderna, har du rätt att arbeta obegränsat under din studietid och du behöver inget särskilt tillstånd för det.
Du kan beviljas uppehållstillstånd i Finland om minst en av dina föräldrar eller mor- eller farföräldrar är eller har varit infödd finsk medborgare.
Om du inte själv är medborgare i ett EU-land, Liechtenstein eller Schweiz men avser att flytta till Finland till en familjemedlem som är EU-medborgare, måste du ansöka om uppehållskort för en familjemedlem till en EU-medborgare.
De flesta kommunerna i Finland är finskspråkiga.
Om du är osäker på om ett visst läkemedel får föras in i Finland ska du fråga råd vid Tullen (Tulli).
En stödbostad kan antingen vara kundens egen ägarbostad, en hyresbostad eller någon annan bostadsform.
Skolan börjar vanligtvis det året då barnet fyller sju år.
Barndagvård och utbildning för barn
Handikappbidrag för vuxna
Vuxnas sexualitetfinska _ svenska _ engelska
Parktanterfinska _ svenska
Vasa
Du behöver inget stort lån för en bostadsrättsbostad.
Många människor får med åldern sämre syn och hörsel.
VAR: Insamlingsställen för farligt avfall, se kierratys.info
Vanligen vårdar någondera av föräldrarna barnet hemma åtminstone under föräldraledigheten (vanhempainvapaa), det vill säga tills barnet är ungefär 9 månader gammalt.
Man kan be om hjälp med sina problem.
hjälpmedelstjänster
linkkiSocial- och hälsovårdsministeriet:
Internationella bortföranden av barnfinska _ svenska _ engelska _ ryska _ franska
Ett hyresavtal kan vara
Rådgivningsbyråns tjänster i den egna kommunen är kostnadsfria.
På rådgivningen får du information om sjukhuset eller sjukhusen i ditt område.
Om begravningsbyråer får du information till exempel från Finlands Begravningsbyråers Förbund (Suomen Hautaustoimistojen Liitto).
Tfn 050 5650 636 (24h)
Antagningsgrunder till yrkesutbildningfinska _ svenska
Du märker väl att vi inte ger råd i hur du ska sköta dina ärenden.
Du får mer information om att leva i Finland med ett handikappat barn på InfoFinlands sida Ett handikappat barn.
Ordna finansiering
Då är föreningen en juridisk person vars medlemmar inte personligen bär ansvar för föreningens verksamhet.
Även utomlands bosatta finska medborgare har rösträtt.
Anbudet kan vara t.ex. 5-10 procent lägre än priset som säljaren har bett om för bostaden.
Dessa aktörer handleder alla som är intresserade av företagande i hela Finland.
Personerna som ska gifta sig ska båda vara närvarande vid vigseln.
Ditt barn kan endast ha ett språk som modersmål.
Information om handikapptjänsternafinska _ svenska _ engelska
ett löneintyg för de senaste sex månaderna före insjuknandet om dina inkomster har ökat.
Arbetspensionsanstalter ordnar yrkesinriktad rehabilitering för arbetstagare.
På utbildningsstyrelsens (Opetushallitus) webbplats finns en sökmotor med vilken du kan kontrollera var och när du kan avlägga examen.
Beviljande av flyktingstatus till asylsökande
För att träffa en hälsovårdare på rådgivningsbyrån för familjeplanering krävs tidsbokning.
Han eller hon ställer dig frågor och bedömer hjälpbehovet.
Helsingfors har goda landsvägsförbindelsermed resten av landet.
Säg upp ditt gamla elavtal innan du flyttar och gör upp ett nytt.
Du kan också fråga direkt av högskolorna.
FPA:s rehabilitering är avsedd för personer som omfattas av den finländska sjukförsäkringen (sairausvakuutus).
Undervisning för invandrare
På InfoFinlands sida Problem i äktenskap och parförhållande finns information om var man kan få hjälp med problem i parförhållanden.
Du kan boka tid vid alla rådgivningsbyråer på samma nummer.
En utredning över grunden för att den person som ansöker om familjeförening vistas i Finland.
Luckan integration
Graviditet och förlossning
Yrkesläroanstalterfinska _ svenska _ engelska
Modersmålsundervisning ges i ryska och i mån av möjlighet även i andra språk.
Förbundet erbjuder även mycket nyttig information och tjänster till synskadade.
Du kan ansöka om en plats
Information om studentexamenfinska _ svenska _ engelska _ franska _ tyska
Utöver detta behöver du en säkerhet för resten av lånesumman.
FPA betalar ut moderskapspenning på samma villkor också till studeranden och arbetslösa.
Finskan har också en del postpositioner.
linkkiInstitutet för de inhemska språken:
Staden ligger i södra Finland vid Finska viken.
Det finns dock fler omständigheter som påverkar den sociala tryggheten, till exempel vilket land du kommer ifrån.
Hur lång boendetid som krävs beror på din situation, vanligtvis ska du ha bott här minst 4–7 år.
Skyddshemmet Mona (turvakoti Mona) är ett skyddshem avsett för invandrarkvinnor och deras barn.
Sådana tjänster är till exempel hälsovård, barndagvård och undervisning.
Om ditt äktenskap slutar med skilsmässa, ändras inte ditt efternamn.
Hindersprövningen görs på magistraten.
Det lönar sig att klä sig varmt eftersom klara nätter vanligtvis också är kalla.
Företagarna i Finland (Suomen Yrittäjät) är företagarnas intressebevakningsorganisation som också producerar sina medlemmar olika tjänster, som till exempel gratis telefonrådgivning i frågor som rör företagande.
Om en asylsökande beviljas flyktingstatus eller uppehållstillstånd på grund av skyddsbehov eller på någon annan grund får han eller hon stanna i Finland.
En make/maka/sambo/partner beviljas inte uppehållstillstånd om förutsättningarna för uppehållstillstånd inte uppfylls.
Då du flyttar till Karleby (Kokkola) ska du registrera dig som invånare i kommunen.
Vid problem hos barn i skolåldern får man hjälp hos skolhälsovårdarna (kouluterveydenhoitaja), skolkuratorerna (koulukuraattori) och socialhandledarna (sosiaaliohjaaja).
Dagvård ordnas också inom familjedagvården och i gruppfamiljedaghem.
Om du vill upprätta ett avtal eller ett testamente för fördelning av egendomen i ett samboförhållande, kan du be om råd till exempel vid rättshjälpsbyrån eller av en jurist.
Ett andelslag är ett företag som ägs av medlemmarna.
Familjedagvård
Rundradion, det vill säga Yle, äger fyra tv-kanaler som visas i hela landet.
Mellersta Österbottens utbildningskoncern erbjuder kurser i finska vid Mellersta Österbottens folkhögskola i Kelviå inom utbildningen i läs- och skrivfärdigheter och den förberedande utbildningen för vuxna invandrare. Det går också att studera finska inom utbildningen som handleder för yrkesutbildning (VALMA) vid Mellersta Österbottens Vuxeninstitut.
linkkiVi läser tillsammans:
Läs mer: Äktenskap.
_ isländska
Myndigheten kan ordna och betala tolkningen när det gäller skötsel av ärenden som behandlas på myndighetens initiativ.
Lämna utrymme runt TV:n, mikrovågsugnen, kylskåpet och frysen.
Tågtrafiken i Finland sköts av bolaget VR.
Nattcaféet finns i Helsingfors på adressen Vasagatan 5, och telefonnumret är 050 443 1068.
Kontaktuppgifter till invandrarenheten:
Var och en får själv välja sin religion.
Kontakta hyresvärden så snart som möjligt och försök förhandla om en förlängning av betalningstiden.
Det kan hända att man i kollektivavtalet har kommit överens om andra villkor och du får lön för en längre tid.
Om du behöver hjälp genast ska du tala om det när du ringer.
Det är snabbt och enkelt att starta företagsverksamhet som enskild näringsidkare.
Tfn 09 2313 9325
Mer information om detta finns på InfoFinlands sida Utländsk examen i Finland.
Om du har tagit ett lån hos en finländsk bank, får skattemyndigheten uppgifterna om lånet direkt från banken.
Om du inte har rätt att använda de offentliga hälsovårdstjänsterna, kan du söka dig till en privat tandläkare.
Mer information hittar du på Vanda stads webbplats.
65101 Vasa
Gator och trafikfinska _ svenska
Ärenden rörande den sociala tryggheten när du flyttar till Finland eller utomlands:
Allemansrätten (jokamiehen oikeudet) är en väsentlig del av den finländska kulturen och lagstiftningen.
För en utvecklingsstörd person är det svårare att lära sig och minnas saker än för andra.
Stöd för närståendevårdfinska
Fråga om verksamheten vid din mödrarådgivning.
Du kan arbeta vid sidan av studierna.
Personförsäkringar kan vara till exempel olycksfallsförsäkring, vårdkostnadsförsäkring och livförsäkring.
Om du behöver besöka tandläkaren snabbt, ta kontakt med social- och hälsostationen i Kilo.
B1 – ASE 3
modersmål
Kvinnan eller mannen kan lämna in skilsmässoansökan på Lapplands tingsrätts kansli i Rovaniemi.
Helsingfors stad betalar dessutom ett kommuntillägg vid hemvårdsstöd till familjer som hemma sköter ett barn som är yngre än två år.
Du kan utnyttja barnrådgivningsbyråns tjänster i din egen kommun om du har hemkommun i Finland.
Rådgivningstjänster hittar du på InfoFinlands sida Ring och fråga om råd.
Du ansöker om stödet från FPA.
Förmedling i familjefrågorfinska _ svenska _ engelska
Du kan också boka tid hos en privatläkare, men kontrollera när du bokar tiden att läkaren har Valviras tillstånd att ge ett utlåtande för abort.
Information om köp av läkemedel hittar du på InfoFinlands sida Läkemedel.
Att hyra en bostadfinska _ svenska _ engelska
Läs mer på InfoFinlands sida Förskoleundervisning.
Elektronisk ansökningsblankett för förskoleundervisningenfinska _ svenska _ engelska
Hälsostationerna har vanligen öppet från måndag till fredag, ungefär kl. 8–16.
Offentliga hälsovårdstjänster
Det öppna universitetet vid Lapplands universitet erbjuder studiemöjligheter enligt studiekraven vid de pedagogiska, juridiska, konst- och samhällsvetenskapliga fakulteterna.
din hemkommun är Vanda
Information för EU-medborgarefinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ rumänska _ ungerska _ italienska
Anställda vid invandrarbyrån
Tänd inte ljus i närheten av till exempel gardinerna, ens om du själv är i rummet.
du inte har för stor förmögenhet.
I Finland finns svenskspråkiga yrkeshögskolor och universitet.
Dessa uppdrag kan vara till exempel:
Du kan hyra ut bostaden till någon annan under högst två år.
På Klockarmalmens begravningsplats finns ett gravområde för konfessionslösa.
Finländska handikapptolkar kan inte nödvändigtvis de teckenspråk som används i andra länder.
Likabehandling
Studiestöd
Tolkningfinska _ engelska
Du kan ringa nödnumret utan riktnummer även om du har ett utländskt mobilabonnemang.
Intyg som utfärdats av en myndighet i ett nordiskt land eller EU-land behöver inte legaliseras.
Om en brand uppstår i din bostad avger brandvarnaren ett högljutt larm och du hinner ut i tid.
Inom dagvården ges även undervisning i finska som andra språk.
linkkiSkatteförvaltningen:
Daghem och andra dagvårdsplatserfinska _ svenska
Barnen undervisas dock inte ännu i läsning.
FPA sköter grundtryggheten i olika skeden av livet för dem som bor i Finland.
Bruksvederlagets storlek beror på bostaden och orten.
InfoFinlands finansiärer har ingått ett samarbetsavtal med vilket man överenskommit om principerna för genomförandet och finansieringen av nättjänsten InfoFinland (tidigare Infobanken) för åren 2017–2020.
Fråga mer vid din egen läroanstalt.
Alla har rätt till integritetsskydd.
Om du blir utvisad, förfaller ditt eventuella giltiga uppehållstillstånd och du måste lämna landet.
Stöd- och serviceboende.
Utmätningsmyndigheten kan även sälja värdefull egendom som du har för att betala skulden.
Asylsökande har inte rätt till finskt socialskydd.
Läs mer: Yrkeshögskolor
Patientombudsmannen ger också information om patientens rättigheter och främjar förverkligandet av dessa.
Du kan få handledning i företagande eller företagarutbildning.
Hyresvärden kan höja hyran i enlighet med vad som anges i hyresavtalet.
Du kan få viktig information om olika organisationers verksamhet och aktuella händelser i olika branscher eller delta i diskussioner.
Om du är arbetslös och söker efter arbete, ska du anmäla dig som arbetssökande hos TE-byrån.
Kurserna i svenska finns under en länk på tjänstens förstasida.
Registreringen är viktig, för utan den kommer du inte att ha rätt till exempelvis social trygghet i Finland.
Dessutom finns det daghem som köptjänst (svenskspråkiga), ett privat daghem och privata familjedagvårdare i Karleby.
Välfärds- och servicepunkten Olkkari
Förskoleundervisningen börjar i augusti.
I Helsingfors finns ett filmarkiv och flera biografer.
Stöd för den blivande modern
Vid magistraten kan du få en finsk personbeteckning, om du inte har ansökt om detta samtidigt som du ansökte om uppehållstillstånd.
Den som vill sluta använda droger kan bli medlem.
Mer information och anmälan finns på NewCo Helsinki webbplats.
Olkkari erbjuder servicehandledning och rådgivning för stadsbor i alla åldrar när det gäller social- och hälsovårdstjänster, kulturella aktiviteter, jobbsökningscoachning, idrottstjänster och organisationsverksamhet.
Torka till exempel inte tvätten ovanför eller i närheten av bastuugnen.
Berätta för hälsovårdaren vilka vaccinationer ditt barn har fått innan ni kom till Finland.
Föräldrarna anmäler sitt barn till förskoleundervisningen vanligtvis i januari eller februari.
Om du planerar att köra bil hem med barnet behöver du ett babyskydd (turvakaukalo) i bilen.
Dessutom är en del av räntan på bostadslånet avdragsgill i beskattningen.
Yles kanaler och flera kommersiella kanaler är avgiftsfria.
Besiktningar görs på besiktningsstationer.
juldagen 25.12
Jourmottagningen vid Haartmanska sjukhuset har öppet vardagar kl. 14–21 och lör–sön kl. 8–21.
I Esbo finns ett vuxengymnasium (aikuislukio) där vuxna kan avlägga gymnasie- och studentexamen.
De första skriftliga källorna om Finland är från 1100–1200-talen. Då anslöts
Intyg om yrkeskunskap med ett fristående yrkesprov
att få veta tidpunkten för intagning för vård om patienten måsta köa till vården
ge arbetstagaren en skriftligt utredning om de centrala villkoren i arbetet
Barnpassningen är avgiftsbelagd.
till skydd utgående från lagar och avtal
linkkiRöda Korset:
Pro-tukipiste har verksamhetsställen i Helsingfors, Tammerfors och Åbo.
Medborgare i ett EU-land, Norge, Island, Lichtenstein och Schweiz kan anmäla sig som arbetssökande via TE-byråns webbtjänst.
I webbtjänsten MinSkatt kan du sköta många skatterelaterade ärenden elektroniskt.
I Karleby finns ungdomsfullmäktige, äldre- och handikappråd samt ett råd för kulturell mångfald.
Civilvigsel äger rum vid magistraten.
Om du flyttar till ett EU-land, ett EES-land eller Schweiz som utsänd arbetstagare (lähetetty työntekijä), ska din arbetsgivare hämta intyget E101/A1 för dig vid Pensionsskyddscentralen.
Integrationstjänster för invandrarefinska _ svenska _ engelska
politiska åsikter.
Du kan ansöka om folkpension om du inte har någon arbetspension eller om din arbetspension är väldigt liten.
du säger upp dig från ditt jobb utan en godtagbar anledning
JA: glasförpackningar (flaskor och matburkar)
Om du har kommit till Finland för att arbeta kan du ha rätt att använda de offentliga hälsovårdstjänsterna i Finland.
Jämlikhet i rekryteringen
Teater och film
Om du har hemkommun i Finland kan du utnyttja de offentliga hälsovårdstjänsterna.
Du hittar kontaktuppgifterna till organisationerna på Handikappforums webbplats.
Information för föräldrar som planerar att skiljasfinska
Ansökan till utbildning
Du kan få finskt medborgarskap
I undantagsfall delas egendomen inte jämnt.
Mer information hittar du vid arbets- och näringsbyrån.
Om du kommer från något annat land till Finland för att studera behöver du en omfattande sjukförsäkring innan du kan få uppehållstillstånd i Finland.
Elektroniskt receptfinska _ svenska _ engelska
Kontaktuppgifter till privata läkare hittar du till exempel på Internet.
Om du kommer från ett EU-land, ett EES-land eller Schweiz till Finland för att studera har du rätt till nödvändig sjukvård med det europeiska sjukvårdskortet.
arbets- och näringsbyrån uppskattar att företagsverksamheten kan vara lönsam
Kontakta rådgivningsbyrån i ditt område genast när du upptäcker att du väntar barn.
Broschyren Information om sexuellt överförda sjukdomar(pdf, 1500kt)finska _ engelska _ ryska _ franska _ somaliska _ arabiska _ kurdiska _ thai
Om arbetstagaren vill att en bedömning av färdigheterna och uppförandet antecknas i arbetsintyget måste arbetsgivaren utfärda ett sådant intyg ännu fem år efter att anställningen har upphört till arbetstagaren på hans eller hennes begäran.
Museer
Läs mer:
Lärare, studiekamrater, bekanta, tidigare kollegor och chefer kan också ingå i ditt nätverk.
Tjänster för företagarefinska _ svenska _ engelska
Fritidsobjekt på kartanfinska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ tyska _ vietnamesiska _ portugisiska _ polska _ holländska _ japanska _ italienska
Observera att du måste legalisera handlingar som har utfärdats av myndigheter utanför EU eller Norden.
Med ett resekort (matkakortti) reser du förmånligare än med kontanter.
Magistraten i Nyland Helsingfors enhet
Om du till exempel avlägger en grundexamen vid universitet, högskola eller yrkeshögskola bör du avlägga 45 studiepoäng under ett läsår för att uppfylla villkoren för fortsatt uppehållstillstånd.
Museerfinska _ svenska _ engelska
Information för hyresgästenfinska _ svenska _ engelska
Brevet innehåller anvisningar om hur du tar emot platsen och hur du anmäler dig.
Detta görs om
Anonyma narkomaner (Nimettömät narkomaanit NA) erbjuder stöd och information samt gruppmöten.
Lekparkerfinska _ svenska _ engelska
du har haft hemkommun i Finland i högst tre år.
Också kyrkans familjerådgivningscentral erbjuder familjerådgivning vid problem i parförhållandet.
Medborgarinstitutetfinska _ svenska _ engelska
Därefter måste du ansöka om uppehållstillstånd eller registrering av EU-medborgares uppehållsrätt för barnet.
FPA och arbetspensionsanstalten bedömer din arbetsförmåga och om du har nytta av rehabilitering.
De kan själva välja hur mycket hjälp som ska ingå i serviceboendet.
Om ditt hem är funktionellt kan du bo hemma även om du har lite svag hälsa.
Du kan även anmäla dig till undervisningen genom att fylla i en blankett, som du får från din egen skola.
Flytta från Finland
Skyddshemmets adress är hemlig.
Social- och hälsovårdsministeriet:
Komihåglistan för dig som flyttar till Finland är avsedd att hjälpa dig med de viktigaste praktiska frågorna som har med flytten att göra.
Gemensam ansökan till gymnasier och yrkesläroanstalterfinska _ svenska
Du kan ansöka till VALMA-utbildningen om du har slutfört grundskolan eller en utbildning som motsvarar grundskolan.
avgångsbetyg från grundskolan med ett godkänt vitsord i finska eller svenska som modersmål eller som andra språk
Vårdbidrag för pensionstagarefinska _ svenska _ engelska
föräldraledighet
Samtal tas emot på följande språk:
Verksamheten är avsedd för alla ungdomar i åldersspannet 13–20 år.
Då kan du avlägga en dubbelexamen (kaksoistutkinto).
partier som finns i partiregistret och
Fler kontaktuppgifter hittar du på Flyktingrådgivningens webbplats.
fälla eller skada växande träd
Blivande förskolebarn får mer information om detta per post, på dagvårdens webbplats och i lokaltidningen.
1550 Helsingfors grundas för att konkurrera med Tallinn om handeln på Östersjön
Läs mer: Stöd- och serviceboende
Då sparas dina personuppgifter, din adress, ditt modersmål och ditt yrke i det finländska befolkningsdatasystemet.
Mer information om hurdana kunskaper de olika nivåerna avser i praktiken får du på Utbildningsstyrelsens (Opetushallitus) webbplats.
linkkiEtuovi.com:
Du kan även låna böcker på bokbussarna.
linkkiFörsvarsmakten:
Arbets- och näringsbyrån (TE-toimisto) ordnar den yrkesinriktade arbetskraftsutbildningen.
Läs mer om gymnasiestudierna på InfoFinlands sida Gymnasium.
Du är själv ansvarig för att skaffa bostad åt dig själv.
Extra kostnader för kläder och matfinska _ svenska
Tolken är antingen på plats eller också kan tolkningen ordnas via telefon eller video.
Företagshälsovården kan dock ge din arbetsgivare en bedömning av huruvida ditt hälsotillstånd tillåter att du fortsätter att arbeta.
I reseplaneraren för cykel- och gångtrafiken kan du söka en lämplig rutt om du vill gå eller cykla.
Synen och hörseln
Den inledande kartläggningen görs vid arbets- och näringsbyrån eller vid kommunen.
Utländskt körkort i Finland
Fpa kan betala grunddagpenning (peruspäiväraha) för en arbetslös företagare som inte är medlem i en arbetslöshetskassa.
Planen kan omfatta t.ex. studier i finska, andra studier eller arbetspraktik.
Familjevård (perhehoito) innebär att en person vårdas, fostras eller omhändertas i ett privat hem utanför det egna hemmet.
Mer information om uppehållstillstånd för studerande och om den sjukförsäkring som krävs för att få uppehållstillstånd får du på Migrationsverkets (Maahanmuuttovirasto) webbplats.
Där kan du vid behov övernatta.
att tvinga någon att sälja sex
Ansökan om uppehållstillstånd för uppstartsföretagare är indelat i två steg:
Om en elapparat börjar brinna, använd inte vatten.
Du kan under utbildningen bekanta dig med olika branscher och fundera på vad du vill studera.
Såväl individer som sambor/gifta par kan ansöka om en hyresetta.
på finska tfn +358 (0)20 692 206
Visa intresse för barnets skolgång och delta till exempel i föräldramöten som skolan ordnar.
Inom forskningen har universitetet två tvärvetenskapliga och internationella
I alla val är det möjligt att rösta också före valdagen, under förhandsröstningstiden.
Positivt beslut
Ett aktiebolag passar för all slags affärsverksamhet.
Läs mer: Tandvård.
intyg på yrkesexamen som du har avlagt på finska eller svenska
Man kan förlora sitt finska medborgarskap om man
I Finland framhävs jämställdhet.
du har fyllt 18 år;
Krishjälp för invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
du har en arbetsplats i Finland och ditt arbetskontrakt är i kraft minst två år
När du vill boka tid för akut tandvård ska du ringa tandvårdens jourtidsbeställning (päivystysajanvaraus) i din hemkommun.
Kamrersvägen 6 A
Du kan söka teaterföreställningar i evenemangskalendrarna på sidorna helsinki.fi och stadissa.fi.
Att framföra vilket som helst motorfordon i onyktert tillstånd (alkohol eller droger) är ett brott.
Läs mer på InfoFinlands sida Bostadslöshet.
För fyrverkerierna har man satt exakta tidsgränser.
Samtidigt som du ansöker om medborgarskap för dig själv, kan du ansöka om det för ett minderårigt barn som du har vårdnaden om.
linkkiUniversitetets almanacksbyrå:
Material från Flerspråkiga bibliotekets samlingar kan lånas från hela Finland.
Kvällstid och under veckoslut har hälsostationen stängt.
undersökningar för att fastställa rehabiliteringsbehovet
Avgiften ska betalas då ansökan ställs.
Du kan också få rätt till den sociala tryggheten i Finland genom att arbeta i Finland.
Också arbetsamhet och flit värdesätts högt.
Fråga mer om kurser i svenska vid din egen arbets- och näringsbyrå.
Om du kommer från ett viseringspliktigt land och ska arbeta i under tre månader, måste du ansöka om ett säsongsarbetsvisum hos den finländska beskickningen.
Uppehållstillståndet kan dock förlängas om du fortsättningsvis har starka band till Finland.
Om du har hemkommun i Finland ska du först kontakta din egen hälsostation (terveysasema).
Även jakt fordrar jakttillstånd.
Klubbarna är avgiftsfria.
Om du har avlagt gymnasiet kan du ansöka till gymnasiebaserad yrkesutbildning (lukiopohjainen ammatillinen koulutus).
Meddela din arbetsgivare om din föräldraledighet två månader innan den börjar.
Läs mer på InfoFinlands sida Behöver du en tolk?
Under våren är vädret ännu svalt, men varmare än på vintern.
Hjälpmedel för arbete och studierfinska _ svenska _ engelska
Vid Stadin ammatti- ja aikuisopisto ordnas förberedande utbildning inför yrkesutbildning för invandrare.
Arbetstagar- och arbetsgivarförbunden förhandlar gemensamt fram branschspecifika kollektivavtal.
Språkstudier i anslutning till annan utbildning
Problemen kan vara till exempel kommunikationssvårigheter, otrogenhet, eller svartsjuka, d.v.s. rädsla för att förlora den andra.
Att lämna Finland
Det erbjuder tjänster för invandrare som bor i Rovaniemi och andra områden i Lapplands län.
Broschyr om besöksförbud(pdf, 418,92 kt)finska _ svenska _ engelska
På 1990-talet ökade inflyttningen från andra länder till Finland.
Fråga om kurserna i finska på din egen arbets- och näringsbyrå.
Byggherrarnas kontaktuppgifterfinska _ svenska _ engelska
fastighetsskatt (kiinteistövero)
Dessutom görs en inledande kartläggning och integrationsplan för invandrare som inte kan registrera sig som arbetslös arbetssökande.
Om skatten inte har betalats, blir du tvungen att betala den i efterskott.
Du måste dock ha ett visum, om du behöver visum till Finland.
studera efter grundläggande studier,
Utöver K.H.Renlunds museum lönar det sig att besöka det naturhistoriska museet Kieppi (Kieppi är stängt tills vidare på grund av brand) samt de många hembygdsmuseerna och övriga de historiska resmålen i regionen.
Dina grannar får inte föra oljud till exempel på nätterna.
Den inkomstrelaterade dagpenningen beräknas utgående från storleken på den lön som du hade innan du blev arbetslös.
I detta fall ska du kontakta magistraten och be om anvisningar om hur barnet registreras.
Tyska
När hälsostationen är stängd, kontakta jourmottagningen på Barnsjukhuset.
Fråga mer vid din egen arbets- och näringsbyrå.
Om du söker asyl i Finland har du rätt till tolkning i ärenden som rör behandlingen av din asylansökan.
linkkiHelsingfors Vuxengymnasium:
Vem som helst kan studera vid ett öppet universitet.
Personer som har sin hemkommun i Esbo har rätt till dessa tjänster.
Tiden räknas från slutet av den månad då du säger upp avtalet.
Läs mer på InfoFinlands sidor Att komma överens om anställningsvillkoren och Innehållet i arbetsavtalet.
Dessutom är det möjligt att ansöka om specialboende, korttidsvård eller tillfällig vård samt handledning hos den öppna vården.
Här menas lagar om social trygghet.)
När en integrationsplan utarbetats kan du få integrationsutbildning.
Om en vara som du köpt har brister ska du först kontakt säljaren.
Läs mer: Ett handikappat barn
Om du har tvingats att sälja sex, kan du även få hjälp vid Pro-tukipiste.
Ni kan komma överens om allt detta på egen hand eller vända er till kommunens socialbyrå (sosiaalitoimisto).
Elektroniska tjänsterfinska _ svenska _ engelska
Då kan du inte söka till en grundskolebaserad yrkesutbildning.
Ekonomihjälp-rådgivningen
Här kan dessutom utländska arbetstagare som ska arbeta i Finland tillfälligt få en finsk personbeteckning utan ett separat besök till magistraten.
Religiös vigsel sker i kyrkan eller ett annat religiöst samfund som har rätt att viga till äktenskap.
I vissa situationer kan tillståndet dock förlängas om du fortfarande har nära anknytning till Finland, till exempel i form av en arbetsplats.
Du kan få grunddagpenning om du omfattas av den sociala tryggheten i Finland utifrån permanent boende eller arbete före arbetslösheten och
När du går hemifrån, kom ihåg att kontrollera att spisen och ugnen och till exempel strykjärnet är avstängda.
Ett tidsbundet avtal innebär att man har avtalat om tidpunkten då arbetet inleds och avslutas.
Undervisning i elevens eget modersmål arrangeras i Karleby på flera olika språk, till exempel under läsåret 2017–2018 arrangerades undervisning på nio olika språk.
Kurser i finska och svenska språket för invandrarefinska
Om du inte har några inkomster, får du föräldradagpenningens minimibelopp.
Du får mer information på InfoFinlands sida Behöver du en tolk?.
Före äktenskapet måste hinder mot äktenskapet prövas.
Om du vill få inkomstrelaterat utkomstskydd för arbetslösa, ska du ansluta dig som medlem i företagarnas arbetslöshetskassa (yrittäjien työttömyyskassa).
linkkiFinlands Simundervisnings- och Livräddningsförbund rf:
Ombudet är en pålitlig vuxen person som hjälper dig med olika ärenden under tiden då Migrationsverket behandlar din ansökan.
Du kan fylla i ansökan på Internet eller posta den till FPA.
Information om arbetarskyddfinska _ svenska _ engelska
Om du behöver mer information om legalisering av handlingar, kontakta magistraten eller utrikesministeriet i ditt hemland.
Högskole- och universitetsutbildningfinska
Man ska göra en anmälan till magistraten när man flyttar till Finland.
Privatföretagare sköter sina premier själva.
På InfoFinlands sida Problem i äktenskap eller parförhållande, får du information om var du kan få råd vid problem i äktenskapet eller i parförhållandet.
Rådgivning på chattenfinska _ svenska _ engelska
Förvalta den bostad vars aktier du äger.
Frivillig återflyttning av flyktingar, asylsökande och emigranter
om du har avlagt studier i ett öppet universitet och söker till ett universitet utifrån dessa studier.
Intressebevakning för företagarefinska _ svenska _ engelska
Var och en får själv välja sin egen religion.
Man försöker emellertid alltid först hjälpa barnet så att det kan bo kvar hemma.
Läkaren kan vid behov skriva remiss till en specialist på gynekologiska polikliniken.
Information om Finland på andra ställen på Internet
Privat tandvård är dyrare än offentlig tandvård.
Märk väl att om räntorna stiger så stiger även lånekostnaderna.
Inkomstregistretfinska _ svenska _ engelska _ ryska _ estniska _ kinesiska
Att få ett skriftligt meddelande i förväg om hyran höjs.
Vid Företagsfinland får du information om olika finansieringsalternativ.
Ofta klarar du dig också på engelska.
Villkor för att du ska få rehabiliterande psykoterapi är att
Skyldighet
Verbböjningengelska
Ett delbeslut av arbets- och näringsbyrån behövs också för tillståndet.
De kan orsaka stora plågor för fåglar och andra djur.
Information om konstundervisningfinska _ engelska
Finländarna är ofta rakt på sak och frispråkighet upplevs inte som något oartigt.
Undervisning för invandrare
Flytta till Finland
Inträdesavgifterna till museerna varierar.
Om du arbetar deltid eller bara lite, bedömer TE-byrån om du kan få en arbetslöshetsförmån samtidigt.
Garantipensionens belopp är mellanskillnaden mellan de övriga pensionerna som du får och garantipensionens fulla belopp.
Huvudstadsregionens skattebyrå betjänar kunderna i centrala Helsingfors.
Om du är under 30 år, kan du fråga råd om jobbsökande på Ohjaamo.
I Vanda finns fyra begravningsplatser som tillhör de evangelisk-lutherska församlingarna.
Om läkemedlet har klassificerats som narkotika är begränsningarna strängare.
Lär dig finska med hjälp av filmerfinska _ engelska _ persiska _ arabiska
Finlands areal är 338 432 km², vilken omfattar landets markområden och insjöar.
Information om klimatet i Finlandfinska _ svenska _ engelska
Religiösa samfund kan hjälpa dig med att ordna begravningen.
Karleby stad betalar extra Karlebystöd för de familjer som tar hand om barn under tre år i hemmet.
Tjänsterna kan vara till exempel hemhjälp, måltidservice, tjänster i anslutning till den personliga hygienen, olika typer av säkerhetstjänster och hälsovårdstjänster.
Om du inte har ingått ett skriftligt uppdragsavtal får bostadsförmedlaren inte kräva dig på förmedlingsarvode.
Läs mer på InfoFinlands sida Rehabilitering.
Dela – kopiera och vidaredistribuera materialet oavsett medium eller format
Du kan ringa skuldlinjen kostnadsfritt från hela Finland och diskutera anonymt dina egna eller en närstående persons ekonomiska bekymmer.
störa hemfriden till exempel genom att slå läger alltför nära en bostad eller genom att föra oväsen
Du måste avtala om utbildningen med TE-byrån innan du inleder utbildningen.
Läs mer: Avfallshantering och återvinning.
Till exempel barnbidrag, moderskapsunderstöd och föräldrapenning betalas även till utlandet.
Gymnasiet tar 2–4 år, beroende på den studerande.
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan man till exempel skapa konst, handarbeten, laga mat, dansa eller idka motion.
Man kan själv be om hjälp hos barnskyddet om föräldrarna är utmattade eller familjen genomgår en svår förändring i livet.
Diskrimineringsombudsmannenfinska _ svenska _ engelska _ ryska _ estniska _ somaliska _ persiska _ arabiska _ kurdiska
Åldringar och handikappade som inte klarar av att bo självständigt, kan bo i ett servicehus eller på en vårdinrättning.
Spara beskattningsbeslutet och den specifikationsdel som du fick på våren tillsammans med skattedeklarationen.
linkkiInstitutet för hälsa och välfärd:
Många länder har en beskickning i Finland.
Information om studentkårer i Finlandfinska _ svenska _ engelska
Om du söker till rehabilitering som ordnas av FPA ska du lämna in din ansökan om rehabilitering till FPA innan rehabiliteringen börjar.
Handpenningen (käsiraha) är en avgift, som betalas för bostaden på förhand.
De högsta statliga organen är riksdagen, presidenten och statsrådet, det vill säga regeringen.
Om föräldrarna inte kommer överens om barnets efternamn, får barnet moderns efternamn.
du inte kan fritt prata om din situation för andra.
Religionens påverkan på arbetslivet
Arbetarskyddsfullmäktige gör sig insatt i arbetarskyddsfrågor som gäller arbetsplatsen, deltar i arbetsplatsens arbetarskyddsinspektioner och informerar de anställda om ärenden som rör arbetets säkerhet och hälsa.
Gå med i InfoFinlands användarpanel här:
Studierna kan även vara tilläggsutbildning eller påbyggnadsutbildning alternativt studier vid universitet eller yrkeshögskola.
Myrbacka hälsostation, Jönsasvägen 4
När ett beslut fattats att ditt boende i Finland är stadigvarande, anses du bo stadigvarande i Finland så länge som
Fråga om kurserna direkt vid vuxengymnasiet.
När hyresavtalet upphör utförs en slutsyn i bostaden.
Också dina tidigare studier kan spela en roll.
Social- och krisjouren (sosiaali- ja kriisipäivystys) hjälper dygnet runt om du eller din familj behöver hjälp i en akut krissituation.
Omatila ordnar vid behov boende för dig och dina barn.
Du kan även bo någon annanstans, men då måste du själv bekosta boendet.
Läs mer: Förlossning.
Det erbjuder tjänster för invandrare som bor i Rovaniemi och andra områden i Lapplands län.
Jag lämnade en ansökan om en kommunal hyresbostad men jag har inte fått en bostad fastän det har gått tid.
Det är oartigt att komma för sent eftersom de andra då tvingas vänta på den som är försenad.
Diskriminering av arbetstagare på grund av deras medlemskap i fackförbund är straffbart.
Studentkåren vid Lapplands universitet informerar också om bostäder som hyrs ut till studerande.
Det är ofta det tryggaste sättet.
I Finland är flaggan något högtidligt.
Ungdomar som oroar sig för sitt eget eller sina föräldrars alkohol- eller drogbruk eller spelande kan kontakta Romppu.
Hur användarna rör sig på webbplatsen
Läs mer på InfoFinlands sida Beskattning.
Du är minst 18 år gammal eller gift.
Stödet betalas inte till utlandet.
Hyresgarantin kan inte användas för att betala hyran för de sista månaderna.
Läs mer: Förlossning
När du ansöker om uppehållstillstånd måste du ha med dig ett pass för att kunna styrka din identitet.
Lagen om jämställdhet mellan kvinnor och män (Tasa-arvolaki) förbjuder diskriminering på grund av kön.
till lön och övriga minimivillkor enligt kollektivavtalet
Föreningar för seniorerfinska _ svenska
InfoFinlands webbplats är responsiv.
Betänketid
Socialbyrånfinska _ svenska
Lapplands universitetfinska _ engelska
Läs mer på InfoFinlands sidor Registrering som invånare.
Bekanta dig med innehållen i InfoFinland före flytten.
Elektroniskt:
Tfn 09 310 44986 (betjänar även på engelska)
Invandrarungdomar kan dessutom studera finska och avlägga grundskolans lärokurs.
Läs mer: Bostadslöshet
Betoningen ligger alltid på den första stavelsen.
I Vanda ordnas yrkesutbildning vid yrkesinstitutet Vantaan ammattiopisto Varia, handelsläroanstalten MERCURIA samt TTS Arbetseffektivitetsföreningen rf:s verksamhetsställe i Vanda.
Där bedrivs det även hobbyklubbar och ordnas kurser och evenemang.
Magisterprogrammet är ett studieprogram som leder till högre högskoleexamen.
Om du inte kommer och inte har avbokat tiden, måste du betala en ersättning.
När du får en studieplats får du rättighet att avlägga båda examina.
Om du behöver brådskande vård, till exempel om du råkar ut för en olycka, har du rätt att genast få vård på jourmottagningen vid den närmaste hälsovårdscentralen eller det närmaste sjukhuset.
Stöd- och serviceboende
Meddela arbetsgivaren om vårdledigheten senast 2 månader innan den börjar.
Ansvar för arbetstagarnas inskolning och säkerhet
Läs mer om språkkunskapskraven på InfoFinlands sida Officiellt intyg över språkkunskaper.
Dagverksamheten kan omfatta till exempel matlagning, motion, samtal och friluftsliv.
Rådgivning för papperslösa utlänningar: 045 2377 104 (måndagar kl. 14–16).
Om du flyttar till Finland för att bo här stadigvarande i minst ett år ska du också registrera dig som invånare i magistraten (maistraatti).
Rehabilitering
Du kan ringa
profilområden: forskning i arktiska och nordliga frågor och forskning inom turism.
linkkiLivsmedelsverket:
Familjen kan anställa en skötare i sitt hem även tillsammans med en annan familj.
Plast (muovi)
Folkhögskolorna (kansanopisto) erbjuder både hobbystudier och yrkesinriktad utbildning.
Du hittar information om skilsmässa på InfoFinlands sida Skilsmässa.
linkkiArbets- och näringsministeriet:
Enligt finländsk lag är en person som är under 18 år ett barn.
I undersökningarna utreds orsaken till barnlösheten.
Om du inte flyttar stadigvarande till Finland, omfattas du vanligen av den sociala tryggheten i Finland så länge din anställning varar.
C1 – ASE 5
Företagarpensionsförsäkringen (FöPL) (YEL-vakuutus) är obligatorisk för företagare i åldern 18–68 år, vars företagsverksamhet inbringar minst 7 799,37 euro om året som arbetsinkomst (år 2019).
Tfn (09) 816 22800
Om du sköter ditt barn hemma kan du delta i Grankulla stads öppna familjeverksamhet. Där kan du träffa andra barnfamiljer.
Du kan söka i den kontinuerliga ansökan även i det fall att du inte fick en studieplats i den gemensamma ansökan.
Fullmäktige väljer ledamöterna till kommunstyrelsen, som har som uppgift att bereda och verkställa fullmäktiges beslut.
Du kan anmäla dig antingen via webbtjänsten eller personligen på TE-byrån.
Du har rätt att arbeta, driva ett företag och studera i Finland med lika villkor som finska medborgare.
Det är bra att komma ihåg att grunden för uppehållstillståndet kan påverka vilka rättigheter du har i Finland.
Som bevis duger till exempel ett utdrag ur boenderegistret eller ett hyreskontrakt med bådas namn.
Du kan rösta i valet till Europaparlamentet om
Österbottens TE-byrå
de grunder enligt vilka lön eller andra vederlag bestäms samt löneperioden
Bibliotek och öppettiderfinska _ svenska _ engelska
Rådgivningen år kostnadsfri.
Första hjälpen-anvisningar för olika situationerfinska _ svenska _ engelska
Människor får ordna möten och demonstrationer och delta i dem.
16 procent har något annat modersmål.
Dagvårdsproducenten måste ha kommunens godkännande.
information om arbetslöshetskassorfinska _ svenska _ engelska
Läs mer: Problem med uppehållstillståndet
Läs också InfoFinlands sida:
Undantag är recept som är utskrivna i de övriga nordiska länderna och europeiska recept. De är giltiga i Finland.
Dessa särskilda tjänster är till exempel färdtjänst, hjälpmedel eller en personlig assistent.
Social trygghet
Kriget slutade med de vitas seger.
Stöd och handledning för unga
Om man är arbetsoförmögen kan man få invalidpension före ålderspensionen.
Information och råd till resenärerfinska _ svenska _ engelska
De finländska myndigheterna intervjuar dessa flyktingar. Utgående från intervjuerna väljer man de flyktingar som tas emot till Finland.
Om du ansöker om en bostadsrättsbostad, behöver du ett ordningsnummer. Du ansöker om ordningsnumret vid Esbo eller Helsingfors stad.
Betala hyran som en girering till hyresvärdens konto.
Om du känner att du behöver information om familjeplanering och prevention kan du kontakta din egen hälsostation.
Telefonnumret till kundrådgivningen och tidsbokningen är (09) 8392 0173.
Ett kollektivavtal kan också vara allmänt bindande.
Fasta hjälpmedel är till exempel stödhandtag, ramper och elektriska dörrar.
Rovaniemi stads välfärds- och servicepunkt ger dig information om stadens tjänster.
Lärarna i årskurserna 7–9 har läst det ämne som de undervisar.
Du kan fiska på Vanda stads fiskeområden i Vanda å, Kervo å och på Finska viken.
kan barnet ges faderns efternamn
Fullmäktigeledamöterna och deras suppleanter väljs vid kommunalval vart fjärde år.
Brottsanmälan kan göras per telefon, personligen på polisstationen eller via polisens webbplats.
Om du vill reservera tid till en läkare ska du ta kontakt med hälsocentralen.
Problem i familjen
Läkemedel från utlandet
Måltidsstöd
Utexaminering från universitetet
Information om svenska språketfinska _ svenska
Du behöver göra så i enlighet med god sed, och inte på ett sätt som ger en bild av att InfoFinland stödjer dig eller ditt användande.
De ungas skyddshus
linkkiViktor Ek:
Flygplatserna i Finlandfinska _ engelska
Varje människa har rätt att delta i samhällslivet.
Regeringen bereder och verkställer riksdagens beslut.
Ta med dig originalexemplaren av de bilagor som krävs för ansökan när du lämnar in din ansökan vid ambassaden eller Migrationsverkets tjänsteställe.
Det räcker med att du anmäler dig.
barnets mor har uppehållsrätt i Finland,
Också i de andra konsthusen i Helsingfors ordnas kulturevenemang för barn och unga.
Om du behöver brådskande vård på kvällen eller veckoslutet, kontakta då jourmottagningen (päivystys).
Du får inte:
På InfoFinlands sida Utbildning i Vanda hittar du information om dagvård för barn i Vanda.
Nätmuseetfinska _ svenska
husdjur
Om du eller din maka/make har hemort i Finland kan du ansöka om skilsmässa enligt Finlands lag.
På sistone har man i läroplanen betonat bland annat helheter som omfattar flera läroämnen, undersökning av vardagliga fenomen samt data- och kommunikationsteknik.
I frågor kring barndagvård och förskoleundervisning kan du också kontakta daghemsföreståndarna eller stadens chef för småbarnsfostran (varhaiskasvatuspäällikkö).
Annan anhörig till en person som fått internationellt skyddfinska _ svenska _ engelska
Mellersta Österbottens yrkesinstitut erbjuder yrkesutbildning i Karleby, Kelviå, Kannus, Kaustby, Perho och Jakobstad.
När du flyttar till Finland
Barn, husdjur eller du själv kan av misstag vrida på spisen.
I många kommuner informerar skolan viktiga ärenden i den webbaserade tjänsten Wilma.
Fråga mer hos din egen samfällighet.
Mer information hittar du på InfoFinlands sida Registrering som invånare.
Ibland kan också personer som inte omfattas av den finländska sjukförsäkringen ha rätt till ersättning från FPA. Fråga mer hos FPA.
Om pengarna inte räcker till för boendekostnaderna fastän du får bostadsbidrag, kan du ansöka om utkomststöd hos FPA.
I Esbo finns också privata tandläkare.
Återkallelse av uppehållstillståndfinska _ svenska _ engelska
Dina möjligheter att få en bostad påverkas av ditt bostadsbehov och dina tillgångar och inkomster.
Webbtjänsten Päihdelinkki
Kontrollera alltid i lönespecifikationen att du har fått rätt belopp.
Du kan tala finska, svenska eller engelska.
Riksdagen (eduskunta) är finska statens viktigaste organ för beslutsfattande.
Planera finansieringen för ditt företag noga innan du grundar företaget.
Om du har rätt till stödet kan du ansöka om stödet hos FPA.
Om du har begått ett brott eller till exempel inte har betalat dina skatter, kan detta utgöra ett hinder för att få finskt medborgarskap.
Institutet erbjuder även undervisning i flera olika språk, bland annat finska, svenska, engelska, tyska, franska, ryska, spanska och italienska.
Grankullavägen 7 02700 Grankulla
Myndigheter såsom daghem eller skola ger information om barnet endast till vårdnadshavaren.
Det underlättar dessutom skötseln av ärenden i banken och med arbetsgivaren.
Språkkaféerfinska _ svenska _ engelska _ ryska
Akademiskt erkännande
Hjälpmedel för hörselnfinska
Om du tar hand om ett under treårigt barn, kan du få hemvårdsstöd (kotihoidon tuki).
Om du gjort ansökningen på internet, kom ihåg att regelbundet kontrollera ditt Enter Finland-konto.
De ordnar verksamhet även för utländska studerande.
att köpa sex av barn under 18 år eller ett offer till människohandel
Dessutom tillhandahåller Flyktingrådgivningen allmän juridisk rådgivning för andra utlänningar.
På rådgivningsbyrån får du anvisningar för en trygg graviditet och förlossning.
Personer under 18 år ska ha minst en vårdnadshavare.
När du uträttar ärenden med statliga myndigheter, till exempel vid arbets- och näringsbyrån (työ- ja elinkeinotoimisto), kan du använda endera språket.
Vi betjänar på finska, engelska, ryska och svenska.
Om du inte flyttar stadigvarande till Finland, kan du i vissa situationer ändå ha rätt att åtminstone delvis omfattas av den sociala tryggheten i Finland medan du arbetar här.
Vissa familjedagvårdare vårdar barnen hemma hos de barn som ingår i gruppen.
Flyttning till eller från Finlandfinska _ svenska _ engelska
Den har format omgivningen i hög grad och bland annat påverkat utvecklingen av hamnverksamheten och handeln.
Skolhälsovården har hand om skolbarns hälsa.
Alla har skyldighet att hjälpa vid en olycka.
att undertrycka och tvinga
I Grankulla finns stadens egna daghem, privata daghem och privata familjedagvårdare.
Om din make/maka/sambo/partner har beviljats asyl eller godkänts som kvotflykting före den 1 juli 2016 och familjen har bildats före hen kom till Finland.
Därefter kan du vid behov kontakta patientombudsmannen (potilasasiamies).
Ansökningen kan tas för behandling först när du besökt beskickningen.
Du ska endast ringa nödcentralen i brådskande nödsituationer, där liv, egendom eller miljön är i fara.
Varje religiöst samfund bestämmer själv vilka villkor vigseln omfattas av och hurdan tillställning vigseln är.
Lånetiden för böckerna är vanligtvis en månad.
I Vanda finns flera läroanstalter som ger grundundervisning i konst speciellt för barn och unga.
Vid högskolorna kan du avlägga högskoleexamen.
Museerna är avsedda för alla.
Polisen anmäler brott som begåtts av barn under 18 år till barnskyddsmyndigheten.
du är asylsökande i Finland och har inte ett giltigt resedokument som berättigar till gränsövergång.
Helsingfors stads rådgivning för invandrare, Helsingfors-info, betjänar alla invandrare i huvudstadsregionen.
Barn till en person som fått internationellt skyddfinska _ svenska _ engelska
Om du vill gå eller cykla i Esbo kan du söka en lämplig rutt i reseplaneraren för cykling och gång.
Företagaren betalar alltså inte skilt ut en lön åt sig.
När en familjemedlem behöver kontinuerlig hjälp och vården är både bindande och krävande, finns det möjlighet att få stöd för närståendevård av kommunen.
Du kan söka till en yrkesinriktad vuxenutbildning om du vill avlägga en examen vid sidan om arbetet.
Om du vill ansöka om ägarbostad i Helsingfors, Esbo eller Vanda, ska du först skaffa ett könummer.
I Finland finns även många läroanstalter som erbjuder studier som inte leder till examen för människor i alla åldrar.
De flesta av FPA:s förmåner är sådana att du har rätt till dem endast om du flyttar ditt stadigvarande boende till Finland.
I ett kompetensbaserat CV kan du gruppera dina färdigheter i olika kompetensområden.
Via den kan du skicka frågor och förslag eller respons till staden.
Faderskapsledigheten får endast tas ut före barnet har fyllt två år.
Den ordnas på våren och hösten.
Om du behöver hjälp med något som rör den mentala hälsan, kan du kontakta mentalvårdsenheten.
Kontrollera ansökningstiden vid den institution där du vill bedriva fortsatta studier.
Karleby blev snabbt en förmögen stad i början av 1800-talet tack vare just handeln med tjära och rederiverksamheten.
Guide om att grunda ett företagfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ turkiska _ kinesiska _ arabiska
Om du har en tillräckligt hög inkomst från arbetet per månad kan du låta din pension vila.
Lapplands studentteaters webbplatsfinska _ engelska
lokal-information
På Migrationsverkets webbplats finns mycket information om uppehållstillstånd.
I Esbo ordnas språkexamina av Axxell och Esbo arbetarinstitut.
Yrkesutbildning som anordnas av arbetsgivaren
Godkännande av reglerna
09 2313 9325 (mån.–fre. kl. 10–12)
Om fett börjar brinna när du lagar mat, kväv elden med till exempel ett kastrullock eller med en släckningsfilt.
du är minst 25 år gammal
På sidan finns information om de situationer då du betraktas ha rätt till den sociala trygghet som grundar sig på boende.
annat identitetsbevis där ditt medborgarskap framgår (om du är medborgare i ett EU-land eller ett nordiskt land)
ett läkarintyg om arbetsoförmögenhet
Stöd under skilsmässan
Om ärendet inte kan lösas på arbetsplatsen, kontakta arbetarskyddsmyndigheterna eller ditt fackförbund.
Rådgivning för invandrarefinska _ engelska _ ryska _ somaliska _ arabiska
På Finnkinos webbplats kan du söka biografer enligt stad på engelska och finska och se vilka filmer som visas.
Information om frågor som rör pensionfinska _ svenska _ engelska _ ryska _ estniska
Gå in på sidan www.infopankki.fi och bekanta dig med Infobankens webbplats.
Kontaktuppgifter till barnatillsyningsmännenfinska _ svenska _ engelska
tekniska områden
Den svenska som talas i Finland kallas finlandssvenska.
Ett tidsbegränsat uppehållstillstånd kan också återkallas om de grunder på vilka tillståndet beviljades inte längre gäller.
En utredning över att du har tillräckliga medel för din försörjning
Diskrimineringsombudsmannen kan ge anvisningar, råd och rekommendationer samt hjälpa med att åstadkomma förlikning i fall som gäller diskriminering.
Också pappor är välkomna till rådgivningen.
Om hälsostationen inte har öppet och situationen är akut, ska du kontakta samjouren vid Pejas sjukhus (Peijaksen sairaalan yhteispäivystys).
Läs mer: Beslutsfattande och påverkan
För utbildningstiden betalas ingen lön.
I Esbo finns många olika föreningar, till exempel kulturföreningar och idrottsklubbar.
Boendekostnaderna varierar mycket.
Vid problem som gäller barn i skolåldern hjälper till exempel skolans hälsovårdare.
Han eller hon kan till exempel inte betala ut en mindre lön än vad som fastställts i kollektivavtalet.
FPA:s och Skatteförvaltningens gemensamma rådgivning hjälper invandrare som har frågor om beskattningen eller den sociala tryggheten.
Skattekortet får du vid skattebyrån.
linkkiVi läser tillsammans-nätverket:
Enheterna för socialt arbete och närarbetefinska _ svenska _ engelska
Farligt avfall (vaarallinen jäte)
intyg på mognadsprov som du har avlagt på finska eller svenska för universitetsexamen eller yrkeshögskoleexamen
Bostaden som du köper täcker en del av säkerheten, vanligen ca 70 procent.
Detta är dock prövningsbaserat, med andra ord är det inte säkert att du får stödet.
Kontaktuppgifter till TE-byråerfinska _ svenska
Att ansöka om kommunal dagvårdfinska _ svenska
Köpa bostad
eller vuxensocialarbetet.
Videoklipp som inte anknyter till tävlingens tema eller är osakliga på andra sätt godkänns inte.
Ge konkreta exempel på ditt kunnande.
Missbruksproblem och spelberoende
skämda och torra livsmedel
Man kan få ersättning först efter att den initiala självrisken (alkuomavastuu) har överskridits, det vill säga efter att du har köpt ersättningsgilla mediciner för över 50 euro under ett år.
TE-byråns tjänster
Återuppbyggnad, industrialisering och kalla kriget 1945–1991
På vissa arbetsplatser kan man köpa förmånliga lunchsedlar som man kan använda på matställen i närheten av arbetsplatsen.
Läkemedelshandel på internetfinska _ svenska _ engelska
Tillräcklig finansiering och noggrann planering är oumbärliga.
Fyll ansökan i tjänsten Studieinfo.fi.
Det ligger bredvid Helsingfors, väster om staden.
Du ansöker om startpenning vid den arbets- och näringsbyrå där du är kund.
Utred i tid när du kan söka.
rätt att resa till Finland och vägra att bli utlämnad till ett annat land
Sexuell hälsa och prevention.
internationalitet (till exempel Europaskolan)
Målet med mödravården är att trygga bästa möjliga hälsa för den gravida modern, fostret, den nyfödda och familjen, förebygga problem under graviditeten och upptäcka dem i ett tidigt skede och vid behov anvisa till fortsatt vård.
Dessutom finns det speciella organisationer för ungdomar, yngre tonåringar och studerande.
Om översättningen görs utomlands måste även översättningen vara legaliserad.
Anställningsrådgivningen har öppet måndag–torsdag klockan 9–11 och 12–15.
För registreringen behöver du ett officiellt identitetskort där ditt medborgarskap framgår eller pass som är i kraft.
På internet finns många bostadsförsäljningsannonser.
Äktenskapsintyget i original (om du är gift)
Insamlingskärl som ofta finns vid husbolaget
Du kan även ansöka om en personbeteckning i Finland vid magistraten eller skattebyrån på din hemort.
Hyrorna för bostäder i Helsingfors grannkommuner (till exempel i Vanda, Esbo eller Kervo) är lite förmånligare än i Helsingfors.
Visste du..?
Du kan även få ersättningen i form av ledighet.
rättshjälpsbyråerna.
Kristelefon på finska: 09 2525 0111
Arbets- och näringsbyråns klienter kan ansöka om arbetslöshetspenning vid FPA.
Information om ortodox vigselfinska _ ryska
Skapa dig ett YouTube-konto och ladda upp videoklippet på YouTube.
Magistraten i Nyland, servicestället i Helsingfors
Till dem hör följande:
Före äktenskap måste man skriftligt begära prövning av äktenskapshinder.
Under moderskapsledigheten får man dock inte arbeta under de två veckor som föregår det beräknade födelsedatumet och under två veckor efter förlossningen.
Därefter tas beslut om tjänsterna, och du kan överklaga beslutet om du inte är nöjd med de tjänster som du har beviljats.
Invandrarmän som har problem med våld kan få hjälp via tjänsten Miehen linja.
Jämlikhet och rättvisa är värden som finländarna skattar högt.
äkta par och registrerade par
Telefonoperatörer i Finlandfinska
Stadigvarande flytt till Finland och stadigvarande boende i Finland
Notera att om du har ett uppehållstillstånd som beviljats på basis av familjeband, så kan förändringar i familjeförhållandena, såsom till exempel skilsmässa, påverka ditt uppehållstillstånd.
Om du önskar kan du ringa förlossningsavdelning då din förlossning satt igång eller om du vill fråga om råd.
Myndigheten betalar dock inte alltid för en tolk.
CV-mallarfinska _ svenska _ engelska _ estniska _ franska _ spanska _ turkiska _ tyska _ portugisiska _ polska _ norska
Yttre religiösa symboler, såsom huvuddukar, är tillåtna i Finland, men de klädregler som gäller på arbetsplatserna måste följas.
Arbetslivet i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ kinesiska _ arabiska
Hälsostationen måste inleda även icke-brådskande vård senast inom tre månader.
Du bör beakta hur uppsägningstiden räknas.
Hjälp till människohandelns offer
Lär mer om mentala tjänster på InfoFinlands sida Mental hälsa.
Studerande från USA kan ansöka om ett Fulbright-stipendium.
linkkiFinlands Dövas Förbund rf:
Du kan fylla i ansökan på Internet, skicka den till FPA per post eller besöka FPA:s kontor.
talförståelse
Tillräckliga medel
Broschyrer om arbetslagstiftningenfinska _ svenska _ engelska
I Finland finns exakta bestämmelser till exempel om hurdant tätskikt ett badrum ska ha.
Det underlättar även skötandet av många officiella ärenden.
Ta kontakt med mödrarådgivningen (äitiysneuvola) i din hemkommun.
Du ser i beskattningsbeslutet om du har betalat rätt mängd skatt.
I vissa fall betalar FPA till exempel ålderspension och familjepension till vissa länder även då du flyttar till landet för över ett år.
Läs mer om bostadsbidrag på InfoFinlands sida Bostadsbidrag.
Läs mer på InfoFinlands sida Finskt medborgarskap.
Om du flyttar till Finland för att arbeta får du vanligtvis rätt till FPA:s förmåner under din anställning, även när din anställning är kortvarig.
Rekreations- och campingområdenfinska _ svenska
Västra Nylands tingsrätt
Ange ditt kontaktspråk till magistraten när du registrerar dig som invånare.
Öppna universitetet (avoin yliopisto) och öppna yrkeshögskolan (avoin ammattikorkeakoulu) ordnar universitets- och yrkeshögskolekurser.
Religionsfriheten för barn och ungafinska
Moninets webbplats
Med hjälp av webbankkoderna kan du till exempel uträtta många myndighetsärenden på nätet.
I Finland gör arbetstagare vanligtvis inte mycket övertid.
Att hyra en bostad
Om du har problem som rör förmedlingsarvodet kan du kontakta Konsumentrådgivningen.
Du kan fråga råd på tjänsten även på nätet genom att fylla i en blankett. Du får svar per e-post.
Tillfälligt boende
Krismottagningen ger dig hjälp och stöd i svåra situationer.
Borgerlig vigsel sker hos magistraten (maistraatti) eller tingsrätten (käräjäoikeus).
Farsdag
Vid födseln, då barnet föds i Finland och faderskapet bekräftas.
Handledd motionfinska _ svenska _ engelska
Du kan anmäla ditt barn till lekparkernas eftermiddagsverksamhet med en anmälningsblankett.
Centret erbjuder bland annat medicinsk undersökning och psykologhjälp.
Om läget är akut, kan du även kontakta social- och krisjouren i Esbo.
Om ni vill ha ett gemensamt efternamn ska ni skicka in en anmälan om namnändring till magistraten.
Hur hittar jag en ägarbostad?
Läs mer: Förskoleundervisning.
Läs mer Den sociala tryggheten i Finland
Då arbetar du kortare dagar och får på motsvarande sätt mindre lön.
Bodelningen kan göras direkt när man har lämnat in den första skilsmässoansökan.
Tfn 029 553 9208
Också i Helsingfors finns det universitet och yrkeshögskolor där man kan studera inom många områden.
Det viktiga är att du har uppehållsrätt i Finland, de yrkeskunskaper som krävs och tillräckliga kunskaper i finska.
Apostilleintyget bevisar att myndighetshandlingen är utfärdad av en behörig person.
Du kan besöka TE-byrån om du inte kan anmäla dig som arbetssökande på nätet eller om du är medborgare i något annat land.
Om du är medborgare i något land som inte tillhör EU och flyttar till Finland som företagare, behöver du antingen ett uppehållstillstånd för företagare, ett uppehållstillstånd för arbetstagare eller ett uppehållstillstånd för uppstartsföretagare.
Talar du engelska/svenska?
Tfn 0295 430291
Kurserna i tjänsten finnishcourses.fi är öppna för alla.
Du måste själv skriftligt begära hindersprövning.
Före äktenskapet måste du begära prövning av äktenskapshinder.
På rådgivningsbyrån följs barnets hälsa och tillväxt.
Klienten får en tid till akutvården, mottagningen eller Min Soite-mottagningen.
Du kan anmäla dig till medborgarinstitutets kurser per telefon eller via internet.
Konsumentrådgivningfinska _ svenska _ engelska
jord- och skogsbruksområden
Vuxengymnasium
Evangelisk-lutherska församlingarfinska
Rättigheter och skyldigheter i en ägarbostad
Åbo
Anmälan till förskottsuppbördsregistret görs med samma anmälan som görs för grundande av företaget, d.v.s. etableringsanmälan (yrityksen perustamisilmoitus).
Kvinnan eller mannen kan lämna skilsmässoansökan i Helsingfors tingsrätts kansli.
Utred din situation tillsammans med socialarbetaren: hur mycket kan du betala i hyra, och kan du få hyresstöd.
En socialarbetare kan hjälpa dig att hitta bostad.
Läs mer: Stöd för vård av barn i hemmet
Mer information finns på Polisens webbplats.
En person kan erhålla flyktingstatus också genom att söka asyl i Finland.
Detta beror på vilken kommun du bor i.
du har bott i Finland i minst fem år med A-tillstånd och
Du kan göra flyttanmälan högst en månad före flyttningsdagen, men den bör göras senast en vecka efter att du har flyttat.
Vid problem i parförhållandet och familjen får man även hjälp av familjerådgivningen vid Vanda församlingar (Vantaan seurakunnan perheneuvonta).
Information om magistraternafinska _ svenska _ engelska
Studierna är inte alltid inriktade på att skaffa ett yrke.
Lapplands arbets- och näringsbyrå
Båda föräldrarna bär ansvaret för underhållet av ett barn under 18 år, även om de inte bor tillsammans.
Vid magistraten (maistraatti) på din egen boningsort kan du ta reda på om du har rätt till en hemkommun i Finland.
Läs mer: Yrkesutbildning.
Information om köp av bostad hittar du på InfoFinlands sida Ägarbostad.
Presentation av e-tjänsten Enter Finland
linkkiExpatFinland.com:
Genomförandet av avtalet följs upp av en styrgrupp.
Hjälp telefonledes
Du kan ansöka om föräldradagpenningar om du omfattas av den sociala tryggheten i Finland och varit sjukförsäkrad i Finland, ett annat EU- eller EES-land eller Schweiz oavbrutet i 180 dagar före det beräknade förslossningsdatumet.
Inte alla företag eller personer som erbjuder hjälp med juridiska ärenden är nödvändigtvis sakkunniga.
Bostad och hemförsäkring
Dolda fel är ofta till exempel fuktproblem.
På InfoFinlands sida När ett barn föds i Finland finns mer information för föräldrar vars barn föds i Finland.
Läs mer om årstiderna i Finland på InfoFinlands sida Klimatet i Finland.
Barnets medborgarskapfinska _ svenska _ engelska
På internet hittar du jobbsajter när du skriver ”avoimet työpaikat” (lediga jobb) i sökmotorns textfält.
Servicerådgivning per telefon
Statsöverhuvud är presidenten, inte en kejsare eller en kung.
Du kan boka tid på hälsostationen per telefon.
Du får ringa nödnumret endast i brådskande nödfall där liv, hälsa, egendom eller miljö är i fara.
InfoFinlands sida Utländska studerande i Finland innehåller viktig information om studielivet i Finland.
är överbefälhavare för Finlands försvarsmakt.
Till samma hushåll hör alla som stadigvarande bor i samma bostad.
De vita fick stöd av Tyskland och de röda av Ryssland.
Lägg till bilagorna alltid i PDF-format.
Seniorinfofinska _ svenska _ engelska
Det finns även stödtjänster i grupp och en möjlighet till umgänge med stöd eller under tillsyn av barnatillsyningsmannen och till sömnskola.
Kondomer kan köpas i butiker, bensinstationer, kiosker och apotek. De kan köpas utan recept.
Yrkesutbildningfinska
14 år
registrering av föreningen.
I Finland värdesätts ärlighet, punktlighet och jämställdhet.
Inkomstrelaterad dagpenning
Du ska ändå lämna in din ansökan i Esbo.
Dickursby hälsostation, Konvaljvägen 11
Fyll i ansökan i tjänsten Opintopolku.fi.
Stöd för närståendevårdfinska _ svenska
Grundläggande information om yrkesutbildningfinska _ svenska _ engelska
Om din hemkommun är tvåspråkig, kan du använda svenska även inom de kommunala tjänsterna, till exempel på hälsostationen.
InfoFinlands webbplats upprätthålls av Helsingfors stad.
Språkkurser
Tjänster för arbetstagare och företagare
linkkiEuropeiska kommissionen:
Ett avtal som bekräftats på detta sätt är lika officiellt som ett domstolsbeslut.
I Finland finns många möjligheter att syssla med musik.
Du kan besöka kliniken utan tidsbeställning torsdagar kl. 14–15.30 eller boka en tid.
En företagare och andra som arbetar åt sig själv kan ordna företagshälsovård för sig själv om de så önskar.
I en förening är det medlemmarna som har makten.
Information om kommunvalfinska _ svenska _ engelska
På den här sidan finns information om tjänsterna i Rovaniemi.
Rådgivning på svenska: 0295 025 510
I Vanda ordnas språkexamina till exempel vid Vanda vuxenutbildningsinstitut (Vantaan aikuisopisto).
Sjukledighet är ingen semester utan den beviljas för att du ska återhämta dig från din sjukdom.
Du får skatteavdrag på samma grunder som andra som bor i Finland stadigvarande.
en minst treårig yrkesinriktad grundexamen
Information för viseringsskyldiga personer
Kurser i finska och svenska språketfinska _ engelska _ ryska
Hemvårdsstödet är skattepliktig inkomst.
Det är i lagen fastställt vilka boendekostnader om kan anses vara skäliga då stödet beräknas.
Vid NewCo Helsinki ordnas informationsmöten om att starta eget för invandrare på finska, engelska, ryska, arabiska och estniska.
Om du ska studera i Finland längre än 90 dagar behöver du ett uppehållstillstånd på grund av studier.
13–21-åriga barn och ungdomar samt deras familjer kan få hjälp hos ungdomscentralen (nuortenkeskus).
Utbildningen kostar alltså inget.
Om du har flyttat till Finland nyligen och behöver stöd med integrationen, kan du få plats i en integrationsutbildning via TE-byrån.
Du kan även lämna panelen när som helst.
Du kan ringa eller skicka e-post.
På InfoFinlands sida Ambassader i Finland hittar du information om andra länders beskickningar i Finland.
Om det inte är möjligt till exempel på grund av barnets läge, fattar läkaren beslut om kejsarsnitt.
Om du kommer till Finland för att arbeta eller som företagare måste du bevisa att ditt arbete eller din företagsverksamhet inbringar dig en tillräcklig utkomst.
Information om storprojekt som förverkligas i regionen och förberedelserna för dessafinska _ engelska _ ryska
Arbets- och näringsbyråer (TE-byråer)
Alla helgons dag är emellertid inte en karneval som Halloween, utan en högtidlig och stilla fest.
Ungefär 7 procent av invånarna är svenskspråkiga och 16 procent har andra modersmål.
På deras webbplatser kan du även ladda ned företagarguider åtminstone på finska och engelska.
Personliga läkemedelfinska _ svenska _ engelska
Vid en tidsbunden anställning kan prövotiden vara högst hälften av den tid anställningen pågår.
Jämställdhetsombudsmannen ger dig även övrig information om lagen om jämställdhet mellan kvinnor och män.
Du måste ansöka separat om denna rätt.
Tjänsterna vid Global Clinic är avgiftsfria för kunderna.
Seniorrådgivningen Tfn: 09 8392 4202
Ansökan om uppehållskort
Om förvaltningsdomstolen avslår besvären kan du i vissa fall ansöka om besvärstillstånd hos högsta förvaltningsdomstolen (korkein hallinto-oikeus).
Den sjunde september 1620 undertecknade Sveriges kung Gustav II Adolf en handling som gav den lilla jordbruks- och fiskebyn vid Ristrand status som stad.
Av plastförpackningar görs nya plastprodukter.
I större städer är det ofta svårare att hitta en lämplig hyresbostad. Även hyran är högre.
allmänt bostadsbidrag
Kroppslig bestraffning av barn är ett brott i Finland.
Om du misstänker att du smittats med en könssjukdom kan du boka tid hos läkaren antingen på hälsostationen eller på en privat läkarstation.
ett land inom Europeiska unionen (EU), ett land inom det Europeiska ekonomiska samarbetsområdet (EES) eller Schweiz eller
Rådgivningarfinska _ svenska
Du kan skicka blanketten per post eller lämna den personligen till magistraten i ditt område.
På varje arbetsplats finns också andra kanaler för den interna kommunikationen, såsom anslagstavlor, e-post eller de anställdas postfack.
Rådgivning till invandrare telefonledes och via e-postfinska _ svenska _ engelska
Polisen inleder utredningen om det finns skäl att misstänka ett brott.
På arbetstid får man inte sköta sina privata angelägenheter, utan detta måste göras utanför arbetstiden.
Familjerådgivningen betjänar barn under 18 år och deras föräldrar.
Om du behöver tolk kan sköterskan på rådgivningsbyrån be en tolk att närvara vid besöken.
I Finland finns några internationella skolor.
Dessa kan vara till exempel arbetslöshetsförsäkring, bostadsbidrag, studiestöd och ekonomiska understöd för barnfamiljer.
Läs mer på InfoFinlands sida Fostran av barn i Finland.
Arbetsgivaren ska se till att jämlikhet och jämställdhet mellan könen förverkligas på arbetsplatsen.
Skilsmässan kan påverka ditt uppehållstillstånd om du har ett tidsbundet uppehållstillstånd på grund av familjeband.
Finland blir självständigt
Du kan söka till en grundskolebaserad yrkesutbildning om du har avlagt lärokursen för den grundläggande utbildningen eller en lärokurs som motsvarar den grundläggande utbildningen.
Radiokanalerna i Finlandfinska
Information om barns och ungas problem finns också på InfoFinlands sida Barns och ungas problem.
Jag avslutade mitt jobb hos min förra arbetsgivare, men jag har inte fått ett arbetsintyg.
Motionsrutter i Karlebyfinska _ svenska
Anmäl alltid förändringar i omständigheterna till FPA.
Medborgarinstituten och arbetarinstituten erbjuder hobbystudier.
På biblioteket kan du låna böcker, tidningar, musik, filmer, spel och mycket annat.
du bott i Finland i minst fyra år med A-tillstånd och
Många finländare pratar bra engelska.
Om du till exempel har en tid klockan tolv, var på plats strax före tolv.
Handikappbidraget beviljas vanligtvis för en bestämd period.
Du kan kontrollera saken vid Fpa.
Under denna tid får du särskild moderskapspenning (erityisäitiysraha).
Vårdnadshavare till en person som fått internationellt skyddfinska _ svenska _ engelska
problem med den mentala hälsan
Staden ordnar tjänster för dem, så att de kan bo självständigt.
Applikationen Suomipassi med flera stödspråkfinska _ engelska
linkkiHelsingfors ortodoxa församling:
Vårdgaranti (hoitotakuu)
Om du också har andra orsaker att vistas i Finland, till exempel en arbetsplats, kan du omfattas av den sociala tryggheten i Finland.
Arbetarskyddsförvaltningen övervakar att de i lagen stadgade arbetarskyddsföreskrifterna följs på arbetsplatserna.
För att kunna studera i ett magisterprogram ska du ha avlagt lägre högskoleexamen.
Du kan inte efteråt kräva ersättning för fel, om
linkkiWordDive:
Utöver detta finns det många museer och museiområden runt omkring i Finland.
För elever som nyligen invandrat finns en klass för förberedande undervisning inför grundskolan vid skolan
Kommunerna kan vara antingen enspråkiga eller tvåspråkiga.
Familjeåterförening
Företagets finansiering kan också delvis bestå av pengar man fått eller lånat. För att ansöka om finansiering ska man ha en ordentlig affärsverksamhetsplan.
Arbetskraftsrådgivare 010 604 6590
Medborgarinstitut och arbetarinstitut
Bondegatan 2
Invandrartjänsterna
Hjälp till offer för familjevåldfinska _ svenska _ engelska
Om du flyttar till Finland av familjeskäl får du vanligen en hemkommun i Finland.
Hjälp till offer för diskriminering
Kommunerna ordnar stödboende och serviceboende för handikappade personer som behöver stöd och hjälp i sitt boende.
I vissa specialfall kan den gälla i fem år.
Arbets- och näringsbyrån
Polisamälanfinska _ svenska _ engelska
Pyhäjoki kommunfinska _ svenska _ engelska
Även en maka/make av samma kön kan få uppehållstillstånd, om ni är gifta eller i ett registrerat parförhållande.
Broschyren HIV i familjen(pdf, 881 kb)finska _ engelska _ ryska
Du kan få personlig rådgivning om startande av ett företag på finska, svenska, engelska, ryska, arabiska, estniska, tyska och italienska.
Barn till en utländsk medborgarefinska _ svenska _ engelska
Du kan avlägga studier vid öppna högskolan fastän du får arbetslöshetsersättning (työttömyyskorvaus).
Om du behöver tillfällig barnpassning i hemmet, kan du kontakta Mannerheims Barnskyddsförbund eller Väestöliitto.
Alla som är bosatta i Finland har rättigheter och skyldigheter enligt lag.
Om du inte har rätt till de offentliga hälsovårdstjänsterna, kan du söka hjälp på en privat läkarstation.
Om du har svårigheter att betala hyran för din bostad ska du ta kontakt med hyresvärden.
I två av gymnasierna i Esbo finns en engelskspråkig IB-linje.
en lämplig yrkeshögskoleexamen eller en annan lämplig högskoleexamen och
Om dina inkomster är små kan du ansöka om bostadsbidrag för bruksvederlaget.
På Grankulla ungdomsgård ordnas många olika slags verksamheter.
Daghem
ökad alkohol- eller droganvändning
Ungdomsbostadsföreningen Rovaniemen nuorisoasunnot ry:s webbplatsfinska
På sidan När ett barn föds i Finland finns viktig information om de praktiska ärenden som du måste ta hand om när barnet har fötts.
Servicestället betjänar invandrare som kommer till Finland för att arbeta i ärenden som berör beskattning och social trygghet.
Du är skyldig
Du avlägger en högre yrkeshögskoleexamen på ungefär ett eller ett och ett halvt år.
Val till Europaparlamentet
Då vårdas akuta sjukdomar och olycksfall på jourmottagningen.
I Finland kan barnen vaccineras (rokotus) mot många smittsamma sjukdomar.
Europeiska sjukvårdskortetfinska _ svenska _ engelska _ estniska _ franska _ spanska _ tyska _ portugisiska _ polska _ holländska _ kroatiska _ rumänska _ ungerska _ italienska
Om ni inte får fram ett avtal där heller, måste ni låta tingsrätten lösa tvisten.
Bibliotekskort
Anmälningar till förskoleundervisningen sker i januari–februari.
Anmälningstiden är vanligtvis i januari.
linkkiKommunförbundet:
Läs mer: Bostadslöshet
Antalet bilagor som krävs till visumansökan kan variera beroende på i vilket land du söker visum.
Ungdomar från Esbo kan också söka till gymnasier i andra städer.
Meddelandet om rösträtt vid ett val skickas hem till dig per post cirka en månad före valdagen.
Intagning för vård måste ske inom sex månader.
Hälsovårdaren följer barnets utveckling, vaccinerar barnet och ger information om rätt kost.
Att begå ett brott har dock påföljder även för personer under 15 år.
För mödrahemmet behöver du en remiss som utfärdas av kommunen.
Hemspråksundervisning för invandrare
De slussar vid behov dig vidare till socialjouren.
Många arbetsgivare använder även Twitter som kommunikationskanal.
På InfoFinlands sida Var hittar jag jobb? hittar du information om jobbsökning i Finland.
På tionde klassen kan du höja dina betyg från grundskolan och du får en plan för fortsatta studier.
Din identitet kan verifieras från en handling som styrker identiteten.
Min tillsvidareanställning upphörde, men min sista lön betalades inte ut.
Flerspråkiga biblioteket ligger i Böle i Helsingfors
Arbetsgivaren får inte betala en lön som är mindre än vad som fastställs i kollektivavtalet.
Brandvarnare säljs i varuhus och järnaffärer.
Som medlem i InfoFinlands användarpanel kan du påverka utvecklingen av webbtjänsten InfoFinland, som finns översatt till flera språk.
Du kan ansöka om plats i den kommunala dagvården via Internet eller med en pappersblankett.
Du kan ansöka om skilsmässa ensam även om din maka eller make inte vill skiljas.
Rättshjälp till flyktingarfinska _ engelska
FPA
Tfn 029 56 61820.
Du kan även ringa och prata på engelska.
Förutsättningar för att få startpeng är bland annat att:
2000 Finland placerar sig på första plats i barns läskunnighet i den första PISA-undersökningen
Läs mer: Mental hälsa
På InfoFinlands sida Hyresbostad får du information om hur du kan hitta en hyresbostad.
Äktenskap och samboförhållande
Ansök om uppehållstillstånd för studerande
I InfoFinland hittar du pålitlig information på ditt eget språk om flytten till Finland, arbetslivet, boende, studier i finska eller svenska språket, utbildning, social trygghet, hälsotjänster, tjänster för familjer, problematiska situationer och fritid.
Jourmottagningen vid
Du kan komma till skyddshemmet dygnet runt.
Även unga kan boka tid hos läkaren och få ett recept för preventivmedel.
linkkiMannerheims Barnskyddsförbund:
Webbtjänsten Infopankki.fi publicerades vid Helsingfors kulturcentral 2003 som ett samarbete mellan Internationella kulturcentret Caisa och Helsingfors stadsbibliotek.
Sjukhusvården räcker vanligen några veckor.
Hjälp med att utarbeta affärsverksamhetsplanen
Finland blev medlem i EU 1995 och var ett av de första länderna som införde euro som valuta.
Många religiösa samfund är verksamma i Vanda och Helsingfors.
Fastlagen
Köpcentret Iso Omena
När du flyttar ut
På InfoFinlands sida Arbeta i Finland hittar du mer information om uppehållstillstånd för arbetstagare.
linkkiÖsterbottens tolkcentral:
Om stöd- eller serviceboende ansöks i hemkommunens socialverk (sosiaalivirasto).
du inte är arbetslös, men går från till exempel lönearbete, studier eller hemmaarbete till företagare
Läs mer på Pensionsskyddscentralens webbplats.
Reservera tillräckliga medel för din försörjning
Den inkomstrelaterade dagpenningen beviljas och utbetalas av den arbetslöshetskassa där du är medlem.
Du kan söka till Finnish for Foreigners-kurserna via öppna universitetet.
Att betala hyran i tid.
Vanligtvis badar man bastu naken.
Personalbranschens regler om rekrytering av utlänningarfinska _ engelska
Modern ska genomgå en läkarundersökning 5–12 veckor efter förlossningen och skicka läkarintyget till FPA.
Om du vill studera i Finland behöver du sannolikt kunna finska.
Utlänningsbyrånfinska _ svenska
För yrkesutbildning förberedande undervisningfinska _ svenska _ engelska
Var kan man beställa en tolk?
Där kan även avlidna som inte är medlemmar i kyrkan begravas.
De får också stöd av förbundets förtroendeman vid konflikter på arbetsplatsen.
Du hittar närmare information om hur du kan söka till en yrkesinriktad vuxenutbildning på InfoFinlands sida Ansökan till utbildning.
Servicehandledningfinska _ svenska
I Finland har alla möjlighet att få kostnadsfri företagsrådgivning.
Om du har uppehållstillstånd och hemkommun i Finland har du rätt att använda de tjänster som kommunen tillhandahåller.
Kontaktuppgifter till vuxensocialarbetetfinska _ svenska _ engelska
Om du vill hitta det förmånligaste priset, kan du jämföra olika elbolags priser.
Dessutom kan nämnden utsätta vite, vilket inskärper förbudet för diskriminering.
Dagvården samarbetar med invandrarbyrån i frågor som rör barnet och familjen.
Separat ansökan
hemma, då familjen anställer en skötare i hemmet
Stadens tjänster för arbetssökande
Sport och motion
Fråga i din hemkommun om förberedande undervisning ordnas på svenska i kommunen.
Karleby polisstation
Väntar du barn ensam eller i en svår livssituation?
Den kan vara baserad på ett jobb, studier, företagsverksamhet, familjeband eller tillräckliga medel.
Information om grundundervisningenfinska _ svenska _ engelska
Bassjälvriskandelens storlek beror på:
Medborgarinstitutetfinska
Somalisktalande klienter 020 634 4905 (mån. och fre. 10–12 och 13–15)
Ta kontakt med handikapprådgivningen som utreder ditt behov av stöd, handledning och tjänster utifrån din situation.
Familjedagvård innebär att skötaren vårdar barnen i sitt eget hem.
Läs mer om att vara arbetsgivare på InfoFinlands sida Arbetsgivarens rättigheter och skyldigheter.
Information om andra möjligheter att studera finska eller svenska hittar du i InfoFinlands avsnitt Finska och svenska språket.
Läs mer: Fritid.
Läs mer på InfoFinlands sida Familjeledigheter.
Santa Sport Spafinska _ engelska
Pulkamontie 6, vån. 2
Asylsökandes uppehållsrätt
Om din vistelse i Finland varar mer än tre månader utan avbrott ska du ansöka om registrering av uppehållsrätten för EU-medborgare i tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
Den grundläggande utbildningen ordnas av kommunerna.
Även korta anställningar eller en praktik kan hjälpa dig att bygga ut ditt nätverk.
Under kvällar och helger är hälsostationerna stängda.
I norra Finland är det mörkare än i södra Finland.
Personen kan dock på grund av sitt handikapp eller sin sjukdom även behöva särskilda tjänster för handikappade för att klara vardagen.
längden på ett tidsbundet arbetsavtal och orsaken till att avtalet är tidsbundet
Då arbetar du kortare dagar och får på motsvarande sätt mindre lön.
MoniNet är ett mångkulturellt center som drivs av Rovalan Setlementti ry och ordnar rådgivning och aktiviteter för invandrare.
Tjänsten är i första hand avsedd för personer med flyktingbakgrund och deras familjemedlemmar.
De offentliga tjänsterna är förmånligare än de privata.
Om du är familjemedlem till en finsk medborgare, behöver din försörjning inte vara tryggad.
Därtill finns det andra stora tätorter i Vanda, till exempel Korso, Björkby-Havukoski, Myrbacka, Mårtensdal, Håkansböle, Västerkulla och Backas.
Om du har ekonomiska problem, lönar det sig för dig att alltid först betala hyran och därefter andra räkningar och skulder.
Trettondagen
Varje arbetsgivare är skyldig att ordna förebyggande företagshälsovård för sina anställda.
Bifoga utlåtandet till din ansökan om uppehållstillstånd för uppstartsföretagare som du skickar till Migrationsverket.
Ordspel för nybörjareengelska _ franska _ japanska
Domstolen tar hänsyn till barnets intressen och dess egna önskemål.
Tjänsten finns på finska och svenska.
Du kan endast söka asyl i Finland på det finska territoriet.
Huvudregeln är att du omfattas av den sociala tryggheten i Finland och har rätt till FPA:s förmåner om du bor stadigvarande i Finland.
Mer information om utbildningsprogram och om ansökan hittar du på läroanstalternas webbplats.
Det är bra att skaffa sig en Internetanslutning så fort som möjligt efter att du har flyttat till Finland.
Om du har en arbetsplats kan din arbetsgivare eventuellt stöda din integration.
Du kan alltså använda samma bibliotekskort på stadsbiblioteken i Vanda, Esbo, Grankulla och Helsingfors.
Om du får ett nekande beslut på din tillståndsansökan kan du överklaga den till förvaltningsdomstolen.
Maken, makan, sambon eller den registrerade partnern till en finsk eller en utländsk medborgare som är bosatt i Finland kan få ett uppehållstillstånd i Finland.
byta lampor
Även en make/maka av samma kön kan få uppehållstillstånd.
Om du behöver råd i frågor kring barns psykiska utveckling, kan du boka en tid hos familjerådgivningen.
Att leva ett normalt liv i ditt hem.
I Helsingfors finns flera grundskolor (peruskoulu).
Familjebandet mellan barnet och föräldern måste bevisas till exempel med en födelseattest med föräldrarnas namn.
Mer information får du på InfoFinlands sida Problem i äktenskap eller parförhållande.
Ansök om dagvårdsplats minst fyra månader innan barnet ska börja i dagvården.
I annat fall måste du betala abonnemanget i förskott.
Legalisering av handlingar
Biograffinska
Om du söker till ett vuxengymnasium, kontakta läroanstalten direkt.
Du kan göra flyttanmälan på internet eller med en blankett som du får i magistraten eller på posten.
Läs mer: Dagvård
Din förälder eller mor- eller farförälder som är beroende av din sambo för sin försörjning
Serviceboende tillhandahålls såväl av kommuner som av privata företag.
Mer information hittar du på föreningens webbplats.
Hemvården omfattar hemtjänster, hemsjukvård och stödtjänster.
Du har rätt att få en inledande kartläggning om
Om du inte har rätt till grunddagpenning eller inkomstrelaterad dagpenning, men omfattas av den sociala tryggheten i Finland, kan du ansöka om arbetsmarknadsstöd.
Mer information får du från ditt hemlands beskickning.
linkkiMoniheli:
Hjälp i hemmet för barnfamiljer(pdf, 500 kb)finska _ engelska
Till klubben ansöker du om plats med samma ansökan om småbarnsfostran (varhaiskasvatushakemus), med vilken du även ansöker om dagvårdsplats.
Ungdomsgårdarfinska
Kommunens hemvård är avgiftsbelagd.
Från NewCo Helsinki får du också hjälp med att utveckla uppstartsföretag.
Du kan granska om du har rätt att arbeta i Finland utan uppehållstillstånd från Migrationsverkets webbplats.
Om du är blind eller har nedsatt syn kan du få tjänster för synskadade.
Identitetskort för utlänningar
I Rovala-institutets utbildning för invandrare kan man studera det finska språket och den finska kulturen, arbetslivsfärdigheter och skaffa sig kunskaper om det finländska samhället.
Yrkesutbildningfinska _ svenska
någon tvingar dig att göra saker som du inte vill göra
Internet- och telefonabonnemangfinska _ svenska _ engelska
Närvarointyg (intyg över att du är studerande vid en läroanstalt som är godkänd i Finland)
Ett nytt efternamn ansöks hos magistraten.
Om du vill kan du även be att en frivillig stödperson som utbildats i att vara stödperson är med på förlossningen.
Registrera ett äktenskap i ditt hemland om du har gift dig i Finland
Migrationsverket ger råd i frågor som rör medborgarskap:
Du kan resa till Finland och de övriga Schengenländerna om du har ett giltigt pass eller något annat resedokument som godkänns i Finland.
Tillsammans med en anställd vid arbets- och näringsbyrån (TE-byrån) gör du en inledande kartläggning och en integrationsplan i samband med att du registrerar dig som arbetssökande.
Handikappade personer kan ha svårt att klara av det dagliga livet på grund av sitt handikapp eller sin sjukdom.
Helsingfors stads webbsidor ger dig information om anmälningsdagen.
Information om Karlebyfinska _ svenska _ engelska
Information om tjänster för barn, ungdomar och familjerfinska _ svenska _ engelska
Du kan ansöka om medborgarskap elektroniskt i tjänsten Enter Finland.
Bifoga din meritförteckning, alltså CV, till ansökan.
Detta innebär att arbetet pågår tills den anställda säger upp sig eller tills arbetsgivaren säger upp den anställda.
Numret till FPA:s pensionsärenden är 020 692 202.
Finland fick flyktingar från många länder och hit flyttade människor med finländskt påbrå från forna Sovjetunionen.
Om du inte har en mekanisk ventilation i ditt hem ska du öppna fönstren och vädra via dem.
Du kan göra en ansökan om föräldradagpenning på FPA:s webbsidor.
Den närmaste flygstationen är Helsingfors–Vanda flygplats.
Om du har frågor om den grundläggande utbildningen kan du kontakta Resultatenheten för den finskspråkiga undervisningen (Suomenkielisen opetuksen tulosyksikkö).
Studentbostäderfinska _ engelska
Du måste i regel själv betala kostnaderna för vården.
Bil och flyg
Läs mer på InfoFinlands sida Nordisk medborgare eller EU-medborgare.
Om du blir utsatt för ett brott
Du kan skaffa könummer i flera olika kommuner.
Tfn (09) 4777 180
Kom till simhallen!(pdf, 2 MB)finska _ svenska _ engelska _ ryska _ estniska _ somaliska _ turkiska _ arabiska _ kurdiska _ thai
Jourmottagningar för barn under 16 år finns i Jorv och på Barnkliniken i Helsingfors.
Även i november och mars kan vädret vara kallt och det kan snöa.
Ett enkel- eller dubbelrum kostar i genomsnitt 60–100 euro per dygn.
Vanligtvis kan inkomstrelaterad dagpenning fås under 400 dagar. Undantag från detta är följande situationer:
Dessutom innehåller InfoFinland länkar till material som publicerats på andra språk.
har barnet rätt att ärva sin far och släkten på sin fars sida och tvärtom
De äldsta av dessa är från 1600-talet.
I Rovaniemi finns 400 bostadsrättsbostäder.
Kyrklig vigsel
Information om den sociala tryggheten i Finlandengelska
Bostadens avfallshantering
Arbetslöshetskassa
Integrationsfrämjande tjänster
Det naturvetenskapliga området
Mer information hittar du på magistratens webbplats.
Du kan personligen registrera dig på Karleby enheten för Magistraten i Västra Finland:
Publicerar och administrerar InfoFinland.
någon hotar med att ange dig till myndigheter om du inte gör som hen säger
Om du ansöker om krävande medicinsk rehabilitering behöver du dessutom en rehabiliteringsplan (kuntoutussuunnitelma).
en yrkesexamen
Du kan avlägga allmän språkexamen i finska eller svenska språket.
Finska medborgare har vissa rättigheter och skyldigheter som utlänningar bosatta i Finland inte nödvändigtvis har.
Du kan få FPA:s studiestöd (opintotuki) om du
Ibland kan begravningen fördröjas på grund av att utredningen av dödsorsaken räcker länge.
Man duar också folk man inte känner, likaså sina kollegor.
Du kan ta reda på biljettpriset på förhand på biografens webbplats.
Ledamöterna till kommunfullmäktige utses i kommunalval som förrättas vart fjärde år.
Det är viktigt att du berättar detta så att hälsovårdaren kan hänvisa dig till öppningsoperation.
Man kommer överens om utförandet av arbetet på gemensamma möten och alla håller fast vid det man kommit överens om.
Boende
Största delen av arbetarinstitutens kurser går på finska eller svenska.
I så fall sköter en av föräldrarna barnet hemma och får en föräldrapenning.
I detta fall räcker det om din sjukförsäkring i första hand täcker läkemedelskostnaderna.
Läs mer: Läkemedel.
På detta inverkar ditt stadigvarande boende och arbete i Finland.
Metall från elapparater (t.ex. guld) återvinns.
Privatpersoner lägger även ut tidningsannonser om bostäder som de hyr ut.
Du kan även gå till Vanda skyddshem (Vantaan turvakoti) eller huvudstadsregionens skyddshem (pääkaupunkiseudun turvakoti).
Stadsborna erbjuds även ett tryggt, omfattande, fungerande och trivsamt nätverk för den lätta trafiken.
Matematik
mån–tors kl. 17–19
Arbetstidsarrangemanget och lönen ska framgå ur avtalet.
Du kan även ansöka om fortsatt uppehållstillstånd på annan grund än för det tidigare tillståndet
Lönen ska vara minst i enlighet med kollektivavtalet eller om inget kollektivavtal finns, uppgå till minst 1211 euro per månad (år 2019).
Om det behövs ytterligare utredningar för din ansökan, kommer detta att meddelas via ditt Enter Finland-konto.
Information på olika språk om mental hälsa på webben
Inom barnskyddet är barnets bästa den högsta prioriteten.
Skyddshemfinska
Metall (metalli)
linkkiUtbildningsstyrelsen:
du är finsk medborgare
Om du begår brott i Finland, kan du även utvisas på grund av brotten.
Om föräldrarna inte är gifta och faderskapet inte har erkänts, är modern barnets vårdnadshavare och bestämmer ensam om alla barnets angelägenheter.
Att se till att även dina gäster följer ordningsreglerna.
Kommunförvaltningenfinska _ svenska _ engelska
Du får inte föra ditt eget avfall till insamlingskärl avsedda för ett annat hus.
När någon som studerat utomlands söker till dessa uppgifter behöver han eller hon oftast Utbildningsstyrelsens avgörande om den tjänstebehörighet som hans eller hennes examen ger.
Utöver dessa finns det flera mindre tätorter, landsbygd och skogar i Esbo.
intyg över lån
FPA betalar ut barnbidrag för varje barn som bor i Finland och omfattas av den sociala tryggheten i Finland.
Beloppet på vattenavgiften beror ofta på det antal personer som bor i bostaden.
Du kan få finskt medborgarskap genom medborgarskapsanmälan (kansalaisuusilmoitus) om du är
Läs mer: Att röra sig i naturen.
förrättar civilvigslar och registrerar parförhållanden,
Råd om jobbsökningfinska _ svenska _ engelska _ spanska
Om din hemkommun är Vanda, kan du få en bostad via Sininauha Oy eller Villenpirtti.
Läs mer på InfoFinlands sidor Bostadsrättsbostad och Delägarbostad.
Stöd till flyktingar
Vid problem som gäller barn under skolåldern, kontakta barnrådgivningen.
Barnet kan även läsa sitt eget modersmål om man har registrerat något annat språk än finska eller svenska som modersmål för barnet.
Tfn (09) 839 23651
I skolan får de unga hjälp av skol- och studenthälsovårdarna (koulu- ja opiskeluterveydenhoitajat), skolkuratorerna (koulukuraattorit) och skolpsykologerna (koulupsykologit).
I hälsovårdstjänsterna vid läroanstalter ordnas också mentalvårdstjänster för studerande.
företagsrådgivning
Om du bor på hyra i ett egnahemshus, ska du ofta betala för uppvärmningen och avfallshanteringen.
En myndig person, alltså en person som har fyllt 18 år, får själv besluta om sin religion.
tfn 020 798 4200
Filmfestivalfinska _ engelska
Vid Esbo bildkonstskola (Espoon kuvataidekoulu) kan barn och unga studera bildkonst.
På Utbildningsstyrelsens webbplats hittar du en förteckning över reglerade yrken och de myndigheter som fattar beslut.
En dag i förskolan
Jämställdhet
Jourmottagningen finns ofta i anslutning till sjukhus, i små städer också i en närliggande stad.
Barnaga, till exempel att slå barnen, är likaså ett brott.
Vid universitet kan man studera i många olika studieområden.
Barnrådgivningen
Tfn (09) 87 100 23
Ring hälsostationen direkt på morgonen när den öppnar.
dina barns födelseattester.
hänga upp en lampa i taket med en upphängningsbygel
Eftermiddagsverksamhetfinska _ engelska
faderns efternamn, om faderskapet har fastställts, eller
I vissa kommunerer separeras inledningsvis biogas från avfallet för att producera el och värme.
Studierna på yrkeshögskola kan vara kostnadsfria eller avgiftsbelagda för studeranden.
sexuellt våld.
Du kan inte inleda din läroavtalsutbildning om du inte har en arbetsplats.
Även barn med funktionsnedsättning kan få tjänster för personer med funktionsnedsättning.
Du får även handledning om hur du sköter ärenden och rådgivning om uppehållstillstånd för arbetstagare.
Arbetslöshetsförsäkring
Egendom
I Vanda finns fem kommunala simhallar.
Problem i parförhållandet
som är infödd finsk medborgare,
Fundera också om du har tillräcklig yrkeskunnighet och erfarenhet och planera hur du ska ordna finansiering.
Telefon: 044 756 7673
bensin
Om du vill kan du samtidigt fortsätta arbeta heltid eller komma överens om en kortare arbetstid med arbetsgivaren.
Längden beror på orsaken till karensen.
I klubben lär sig barnet tala finska, fungera i en grupp och där kan barnet träffa andra barn.
Flykting
Kurser för invandrarefinska _ engelska _ ryska
Om inte hinner studera finska vid din egen läroanstalt, finns det kurser i finska vid många andra läroanstalter.
Kyrklig vigsel kan förrättas i
Verksamheten av Mellersta Österbottens Nyföretagarcentral FIRMAXI fortsätter som en del av KOSEKs tjänster.
Öppningsoperationen gör förlossningen och undersökningarna under graviditeten lättare.
Betalningsanmärkning
Ansökan för examensstuderande
ELY-centralernafinska _ svenska _ engelska
I Finland finns även många allmännyttiga samfund som har förmånliga hyresbostäder.
inte uppfyller arbetsvillkoret, d.v.s. inte arbetat tillräckligt länge innan du blev arbetslös eller fått förvärvsrelaterad dagpenning eller grunddagpenning under maximitiden.
Ring nödnumret endast om det handlar om ett nödfall, till exempel en akut sjukdomsattack.
Du får inte arbeta på en byggplats utan namnskylt.
Om du studerar vid en högskola får du också måltidsstöd (ateriatuki).
Om du har uppehållstillstånd på grund av familjeband, har du rätt att arbeta och studera i Finland.
Du kan söka till en yrkesinriktad vuxenutbildning också om du har avlagt en yrkesexamen eller en högskoleexamen.
Boende i bostadsrättsbostad
Vid Esbo arbetarinstitut (Espoon työväenopisto) kan du studera till exempel språk, handarbete och matlagning eller delta i ledd motion.
Ingen kan heller mot sin vilja tvingas att delta i religionsutövande.
Om du inte kan göra ansökan på internet eller inte vet hur man gör det kan du också lämna in en pappersansökan jämte bilagor vid Finlands beskickning närmast dig.
Via dessa sidor hittar du snabbt den information som du behöver i kortfattade form.
Information om tuberkulosfinska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Vid Centria yrkeshögskola kan man avlägga högskoleexamen i teknik, företagsekonomi, social- och hälsovård.
Hälsomotion för personer i arbetsför ålderfinska
viktiga affärsförhandlingar som pågår längre än väntat.
Tfn 040 489 2129
Antagning enligt prövningfinska _ svenska
nivåerna C1 och C2: en avancerad språkanvändares språkkunskaper (taitavan kielenkäyttäjän kielitaito)
Utbildningen är avsedd för unga som vill studera på gymnasiet, men vars språkkunskaper inte är tillräckliga för gymnasiestudier.
Receptet skrivs ut av en läkare.
Handlingen ska vara legaliserad för att magistraten ska kunna föra in dina uppgifter i befolkningsdatasystemet.
Anteckna allt detta i din affärsverksamhetsplan.
Om du vill komma till Finland som utbytesstudent ska du kontakta till exempel studentexpeditionen eller den internationella enheten vid din egen läroanstalt.
Den uttalas lite annorlunda än den svenska som talas i Sverige.
Barnets andra förälder kan vara med på förlossningen.
Man kan inte köpa en bostadsrättsbostad.
Närmare uppgifter om integrationsplanen finns på InfoFinlands sida Integration i Finland.
Frivillig utbildning med arbetslöshetsförmån
Utöver en ersättning kan kommunen ordna även andra tjänster genom vilka vården i hemmet stöds.
Väestöliitto erbjuder parrådgivning och parterapi på finska och engelska.
I vissa fall kan du dock bibehålla din rätt till den sociala tryggheten i Finland även om du vistas utomlands över ett år.
Finland tar som kvotflyktingar emot personer som har flyktingstatus enligt
Barn och unga kan delta i grundläggande undervisning i musik, dans, bildkonst och hantverk.
Om du har rätt till moderskapsunderstöd, moderskapspenning eller andra understöd, ska du ansöka om dem vid FPA.
Om du får ett uppehållstillstånd i Finland registreras du automatiskt i det finska befolkningsdatasystemet.
Läs mer om avgifterna för en hyresbostad, till exempel hyresdeposition, på InfoFinlands sida Hyresavtal.
disponering av barnets egendom
Också utlänningar, d.v.s. personer som inte har finskt medborgarskap, kan grunda en registrerad förening.
Idrottsklubbarfinska _ svenska _ engelska
I Esbo finns flera tåg- och metrostationer.
Religiösa grupper måste inte registrera sig som samfund, utan de kan även verka utan att ha registrerat sig.
Asylsökande har inte rätt till familjeåterförening.
I Esbo finns elva finskspråkiga och ett svenskspråkigt gymnasium (lukio).
Öppettiderna för Lapplands TE-byrå
Hos en privat hyresvärd kan det gå snabbt att få en bostad, men hyran kan vara högre än i stadens hyresbostäder.
Registrering av utlänningarfinska _ svenska _ engelska
Broschyr om erkännande av examen(pdf, 102,14 kt)finska _ svenska _ engelska _ ryska _ estniska _ franska _ spanska _ kinesiska _ persiska _ arabiska _ portugisiska
Tips för boende(pdf, 1,5 Mt)finska _ engelska _ ryska _ somaliska _ arabiska _ kurdiska
Ansök om uppehållstillstånd för uppstartsföretagare och besök Finlands beskickning eller Migrationsverkets serviceställe för att styrka din identitet.
Godkända läroanstalter är läroanstalter efter grundskolan, till exempel universitet, högskolor och yrkesläroanstalter.
Rovaniemi yrkeshögskola eller RAMK är den nordligaste yrkeshögskolan inom EU. Skolan ingår i Lapplands högskolekoncern.
Stödets storlek och villkoren för att erhålla stödet kan variera mellan olika kommuner.
Konsumentskyddslagen tryggar konsumentens rättigheter i Finland.
TE-byrån gör den inledande kartläggningen.
Om du har rätt till arbetslöshetsersättning i ditt hemland, kan du även få den tillfälligt utbetald till Finland.
Rovaniemi yrkeshögskola
Stöd för privat vårdfinska _ svenska _ engelska
Det är inte ovanligt att söka hjälp för att få stöd med den mentala hälsan.
Du kan vara med i invånarverksamheten eller ta ett invånarinitiativ.
Om arbetet upphör och arbetstagaren blir arbetslös kan han eller hon ansöka om inkomstrelaterad arbetslöshetsdagpenning från kassan.
Helsingfors har cirka 600 000 invånare. 83 procent av invånarna har finska och 6 procent har svenska som modersmål.
Du måste ansöka om plats i förskoleundervisningen.
Om du har frågor kring fordonsskatten eller anmälan om ibruktagande, kan du ringa skatteförvaltningens telefontjänst:
Du kan inte få ett kontinuerligt tillstånd på basis av studier.
I Vanda finns även en internationell skola, där man kan avlägga grundskolan på engelska.
Organisationssmedjanfinska _ svenska _ engelska
Mervärdesskatt
Information om fackförbundsverksamhetfinska _ svenska _ engelska _ ryska _ estniska _ franska
Om du är EU-medborgare kan du ansöka om permanent uppehållsrätt när du har bott i Finland fem år.
Lämna inte brinnande ljus utan uppsikt.
Nyföretagarcentraler
Esbo stads rådgivning för seniorer
Rådgivningstjänster
Arbetskraftsutbildningen är avsedd för arbetslösa arbetssökande.
Lyft fram sådant som är viktigt i arbetsuppgiften.
Om dina studier i Finland pågår högst tre månader behöver du inget uppehållstillstånd.
När hälsostationen har stängt ska du kontakta jourmottagningen vid Barnsjukhuset.
Felaktigt ifyllda ansökningar tas inte emot.
Underhållsbidraget är ett bidrag som den förälder som inte bor med barnet betalar för att delta i barnets levnadskostnader.
Om du är medborgare i ett EU-land, får du sannolikt inte asyl i Finland.
Alla får själva välja sin bostadsort och röra sig fritt i Finland.
linkkiYle.fi:
linkkiIESAF:
