Då upphörde Saul att förfölja David och drog mot filistéerna. Därav fick det stället namnet Sela-Hammalekot.
Men själva kunna vi icke åt dem giva hustrur av våra döttrar, ty Israels barn hava svurit och sagt: Förbannad vare den som giver en hustru åt Benjamin.»
Då gingo de fem männen vidare och kommo till Lais; och de sågo huru folket därinne bodde i trygghet, på sidoniernas sätt, stilla och trygga, och att ingen gjorde någon skada i landet genom att tillvälla sig makten; och de bodde långt ifrån sidonierna och hade intet att skaffa med andra människor.
Filippus skyndade fram och hörde att han läste profeten Esaias. Då frågade han: »Förstår du vad du läser?»
jag vill lyfta mina händer upp till dina bud, ty de äro mig kära, och jag vill begrunda dina stadgar.
De omringa mig, ja, de omringa mig, men i HERRENS namn skall jag förgöra dem.
Och var och en av dem förde med sig skänker: föremål av silver och av guld, kläder, vapen, välluktande kryddor, hästar och mulåsnor. Så skedde år efter år.
då berövas de ogudaktiga sitt ljus, och den arm som lyftes för högt brytes sönder.
Den rättfärdiges förvärv bliver honom till liv; den ogudaktiges vinning bliver honom till synd.
Men Jojada blev gammal och mätt på att leva och dog så; ett hundra trettio år gammal var han vid sin död.
Och de gjorde så och läto dem alla lägga sig ned.
Och när de så, under sin flykt för Israel, hade kommit till den sluttning som går ned från Bet-Horon, lät HERREN stora stenar falla över dem från himmelen, hela vägen ända till Aseka, så att de blevo dödade; de som dödades genom hagelstenarna voro till och med flera än de som Israels barn dräpte med svärd.
Och Jesus växte till i ålder och vishet och nåd inför Gud och människor.
Och det fick en mun sig given, som talade stora ord och vad hädiskt var, och det fick makt att så göra under fyrtiotvå månader.
de skulle nämligen fråga prästerna i HERREN Sebaots hus och profeterna sålunda: »Skola vi framgent hålla gråtodag och späka oss i femte månaden, såsom vi hava gjort nu i så många år?»
den fostrar oss till att avsäga oss all ogudaktighet och alla världsliga begärelser, och till att leva tuktigt och rättfärdigt och gudfruktigt i den tidsålder som nu är,
Och konungen ropade med hög röst och befallde att man skulle hämta besvärjarna, kaldéerna ock stjärntydarna. Och konungen lät säga så till de vise i Babel: »Vemhelst som kan läsa denna skrift och meddela mig dess uttydning, han skall bliva klädd i purpur, och den gyllene kedjan skall hängas om hans hals, och han skall bliva den tredje herren i riket.»
Och när man hade offrat brännoffret, sade Jehu till drabanterna och kämparna: »Gån in och slån ned dem; låten ingen komma ut.» Och de slogo dem med svärdsegg, och drabanterna och kämparna kastade undan deras kroppar. Därefter gingo de in i det inre av Baals tempel
Och det skall ske på den tiden att jag skall göra Jerusalem till en lyftesten för alla folk; var och en som försöker lyfta den skall illa sarga sig därpå. Och alla jordens folk skola församla sig mot det.
Och prästen skall av offret taga en handfull, det som utgör själva altaroffret, och förbränna det på altaret; därefter skall han giva kvinnan vattnet att dricka.
Hälsen alla bröderna med en helig kyss.
vidare Ajalon med dess utmarker och Gat-Rimmon med dess utmarker;
Och ändå säga de av Israels hus: »Herrens väg är icke alltid densamma»! Skulle verkligen mina vägar icke alltid vara desamma, I av Israels hus? Är det icke fastmer eder väg som icke alltid är densamma?
Men kommen ihåg, I mina älskade, vad som har blivit förutsagt av vår Herres, Jesu Kristi, apostlar,
Till de andra åter säger jag själv, icke Herren: Om någon som hör till bröderna har en hustru som icke är troende, och denna är villig att leva tillsammans med honom, så må han icke förskjuta henne.
Vi vilja icke lämna eder, käre bröder, i okunnighet om huru det förhåller sig med dem som avsomna, för att I icke skolen sörja såsom de andra, de som icke hava något hopp.
Och i första månaden, på fjortonde dagen i månaden, är HERRENS påsk.
är en man som bedrager sin nästa och sedan säger: »Jag gjorde det ju på skämt.»
Nej, hellre vill jag nu bliva kvävd, hellre dö än vara blott knotor!
Han som icke har skonat sin egen Son, utan utgivit honom för oss alla, huru skulle han kunna annat än också skänka oss allt med honom?
Så skall det gå den glada staden, som satt så trygg, och som sade i sitt hjärta: »Jag och ingen annan!» Huru har den icke blivit en ödemark, en lägerstad för vilda djur! Alla som gå där fram skola vissla åt den och slå ihop händerna.
Såsom HERREN hade bjudit Mose så hade Israels barn i alla stycken gjort allt arbete.
de hava öron och lyssna icke till, och ingen ande är i deras mun.
Med honom är en arm av kött, men med oss är HERREN, vår Gud, och han skall hjälpa oss och föra våra krig. Och folket tryggade sig vid Hiskias, Juda konungs, ord.
Men det skall ske att var och en som åkallar HERRENS namn han skall varda frälst. Ty på Sions berg och i Jerusalem skall finnas en räddad skara, såsom HERREN har sagt; och till de undsluppna skola höra de som HERREN kallar.
Då räckte Aron ut sin hand över Egyptens vatten, och paddor stego upp och övertäckte Egyptens land.
Så gick Åklagaren bort ifrån HERRENS ansikte och slog Job med svåra bulnader, ifrån fotbladet ända till hjässan.
Och jag betraktade det och gav akt därpå; då fick jag däri se fyrfota djur, sådana som leva på jorden, tama och vilda, så ock krälande djur och himmelens fåglar.
En annan sträcka sattes i stånd av Malkia, Harims son, och av Hassub, Pahat-Moabs son, och därjämte Ugnstornet.
Därefter sade han: »Tag pilarna.» Och när han hade tagit dem, sade han till Israels konung: »Slå på jorden.» Då slog han tre gånger och sedan höll han upp.
Femton alnar högt steg vattnet över bergen, så att de övertäcktes.
I två hela år bodde han sedan kvar i en bostad som han själv hade hyrt. Och alla som kommo till honom tog han emot;
Hos honom är väldighet och förskräckande makt, hos honom, som skapar frid i sina himlars höjd.
Och därvid kommer det icke an på om någon är grek eller jude, omskuren eller oomskuren, barbar eller skyt, träl eller fri; nej, Kristus är allt och i alla.
Sedan gick allt folket hem, var och en till sitt; men David vände om för att hälsa sitt husfolk.
Sina gärningars kraft har han gjort kunnig för sitt folk, i det han gav dem hedningarnas arvedel.
Och han skall döma mellan hednafolken och skipa rätt åt många folk. Då skola de smida sina svärd till plogbillar och sina spjut till vingårdsknivar. Folken skola ej mer lyfta svärd mot varandra och icke mer lära sig att strida.
fursten Dison, fursten Eser, fursten Disan. Dessa voro horéernas stamfurstar i Seirs land, var furste för sig.
När jag vill hela Israel, då uppenbarar sig Efraims missgärning och Samariens ondska. Ty de öva falskhet, tjuvar göra inbrott, rövarskaror plundra på vägarna.
Och Israel kom till Egypten, Jakob blev en gäst i Hams land.
Då alltså Edom icke tillstadde Israel att tåga genom sitt område, vek Israel av och gick undan för honom.
Onda andar blevo ock utdrivna ur många, och de ropade därvid och sade: »Du är Guds Son.» Men han tilltalade dem strängt och tillsade dem att icke säga något, eftersom de visste att han var Messias.
Ty jag är HERREN, som har fört eder upp ur Egyptens land, för att jag skall vara eder Gud. Så skolen I nu vara heliga, ty jag är helig.
Och jag skall sätta dem till att förrätta tjänsten i huset vid allt tjänararbete där, allt som där skall utföras.
av fäkreatur sjuttiotvå tusen,
Begär av mig, så skall jag giva dig hedningarna till arvedel och jordens ändar till egendom.
Om någon icke förbliver i mig, så kastas han ut såsom en avbruten gren och förtorkas; och man samlar tillhopa sådana grenar och kastar dem i elden, och de brännas upp.
Och städerna Sodom och Gomorra lade han i aska och dömde dem till att omstörtas; han gjorde dem så till ett varnande exempel för kommande tiders ogudaktiga människor.
Då han nu vandrade utmed Galileiska sjön, fick han se två bröder, Simon, som kallas Petrus, och Andreas, hans broder, kasta ut nät i sjön, ty de voro fiskare.
Sannerligen säger jag eder: Den stund kommer, jag, den är redan inne, så de döda skola höra Guds Sons röst, och de som höra den skola bliva levande.
Var och en som hatar sin broder, han är en mandråpare; och I veten att ingen mandråpare har evigt liv förblivande i sig.
Men i stället hängåven I eder åt fröjd och glädje; I dödaden oxar och slaktaden får, I åten kött och drucken vin, I saden: »Låtom oss äta och dricka, ty i morgon måste vi dö.»
Och vilddjuret, som jag såg, liknade en panter, men det hade fötter såsom en björn och gap såsom ett lejon. Och draken gav det sin makt och sin tron och gav det stor myndighet.
i andra raden en karbunkel, en safir och en kalcedon;
Om du stötte den oförnuftige mortel med en stöt, bland grynen, så skulle hans oförnuft ändå gå ur honom.
Och det vart afton, och det vart morgon, den femte dagen.
Och denna stadga skall du hålla på bestämd tid, år efter år.
Sedan de hade ätit sig mätta, lättade de skeppet genom att kasta vetelasten i havet.
Detta blev en orsak till synd; folket gick ända till Dan för att träda fram inför den ena av dem.
HERREN är rättfärdig därinne, han gör intet orätt. var morgon låter han sin rätt gå fram i ljuset, den utebliver aldrig; men de orättfärdiga veta icke av någon skam.
Om du ser att den fattige förtryckes, och att rätt och rättfärdighet våldföres i landet, så förundra dig icke däröver; ty på den höge vaktar en högre, och andra ännu högre vakta på dem båda.
Noa, Sem, Ham och Jafet.
Se, detta står upptecknat inför mina ögon; jag skall icke tiga, förrän jag har givit vedergällning, ja, vedergällning i deras sköte,
Alltså, att han som förlänade eder Anden och utförde kraftgärningar bland eder gjorde detta, kom det sig av laggärningar eller därav att I lyssnaden i tro,
Men hennes handelsförvärv och vad hon får såsom skökolön skall vara helgat åt HERREN; det skall icke läggas upp och icke gömmas, utan de som bo inför HERRENS ansikte skola av hennes handelsförvärv hava mat till fyllest och präktiga kläder.
I den församling som fanns i Antiokia verkade nu såsom profeter och lärare Barnabas och Simeon, som kallades Niger, och Lucius från Cyrene, så ock Manaen, landsfursten Herodes' fosterbroder, och Saulus.
Ty HERREN Gud är sol och sköld; HERREN giver nåd och ära; han vägrar icke dem något gott, som vandra i ostrafflighet.
Se, dagar skola komma, säger HERREN, då jag skall låta en rättfärdig telning uppstå åt David. Han skall regera såsom konung och hava framgång, och han skall skaffa rätt och rättfärdighet på jorden.
Då bugade sig Bat-Seba, med ansiktet mot jorden, och föll ned för konungen och sade: »Må min herre, konung David, leva evinnerligen!»
Och jag skall göra dem till ett enda folk i landet, på Israels berg; en och samma konung skola de alla hava; de skola icke mer vara två folk och icke mer vara delade i två riken.
För kehatiternas släkter föll lotten ut så, att bland dessa leviter prästen Arons söner genom lotten fingo ur Juda stam, ur simeoniternas stam och ur Benjamins stam tretton städer.
Och alla flyktingar ur alla hans härskaror skola falla för svärd, och om några bliva räddade, så skola de varda förströdda åt alla väderstreck. Och I skolen förnimma att jag, HERREN, har talat.
Ty konungen hade en egen Tarsisflotta på havet jämte Hirams flotta; en gång vart tredje år kom Tarsisflottan hem och förde med sig guld och silver, elfenben, apor och påfåglar.
Låt min muns frivilliga offer behaga dig, HERRE, och lär mig dina rätter.
Det ena som det andra har jag sett under mina fåfängliga dagar: mången rättfärdig som har förgåtts i sin rättfärdighet, och mången orättfärdig som länge har fått leva i sin ondska.
Dock, huru skulle det kunna få ro, då det är HERRENS bud det utför? Mot Askelon, mot Kustlandet vid havet, mot dem har han bestämt det.
Då sade han till sina tjänare: »I sen att Joab där har ett åkerstycke vid sidan av mitt, och på det har han korn; gån nu dit och tänden eld därpå.» Så tände då Absaloms tjänare eld på åkerstycket.
Och närmast Simeons område skall Isaskar hava en lott, från östra sidan till västra.
Och Saul talade med sin son Jonatan och med alla sina tjänare om att döda David; men Sauls son Jonatan var David mycket tillgiven.
Den som tror och bliver döpt, han skall bliva frälst; men den som icke tror, han skall bliva fördömd.
och min ande fröjdar sig i Gud, min Frälsare.
Så äro vi då alltid vid gott mod. Vi veta väl att vi äro borta ifrån Herren, så länge vi äro hemma i kroppen;
Då gick han åstad och begynte förkunna i Dekapolis huru stora ting Jesus hade gjort med honom; och alla förundrade sig.
Och hela Juda gladde sig över eden; ty de hade svurit den av allt sitt hjärta, och de sökte HERREN med hela sin vilja, och han lät sig finnas av dem, och han lät dem få ro på alla sidor.
så må du veta: när profeten talar i HERRENS namn, och det som han har talat icke sker och icke inträffar, då är detta något som HERREN icke har talat; i förmätenhet har då profeten talat det; du skall icke frukta för honom.»
Sedan fick jag i min syn höra en örn, som flög fram uppe i himlarymden, ropa med hög röst: »Ve, ve, ve över jordens inbyggare, när de tre övriga änglar, som skola stöta i basun, låta sina basuner ljuda!»
Jag skyndar mig och dröjer icke att hålla dina bud.
Hos dig må icke finnas någon som låter sin son eller dotter gå genom eld, eller som befattar sig med trolldom eller teckentydning eller svartkonst eller häxeri,
Och varen framför allt uthålliga i eder kärlek till varandra, ty »kärleken överskyler en myckenhet av synder».
Och såsom han uttydde för oss, så gick det. Jag blev åter insatt på min plats, och den andre blev upphängd.»
Såsom ditt namn, o Gud, så når ock ditt lov intill jordens ändar; din högra hand är full av rättfärdighet.
Och må nu icke mitt blod falla på jorden fjärran ifrån HERRENS ansikte, då Israels konung har dragit ut för att söka efter en enda liten loppa, såsom man jagar rapphöns på bergen.»
Av invånarna i Bet-Semes blevo ock många slagna, därför att de hade sett på HERRENS ark; han slog sjuttio man bland folket, femtio tusen man. Och folket sörjde däröver att HERREN hade slagit så många bland folket.
Han kan icke undslippa mörkret; hans telningar skola förtorka av hetta, och själv skall han förgås genom Guds muns anda.
Och detta är lagen om spisoffret: Arons söner skola bära fram det inför HERRENS ansikte, till altaret.
och sade: »Om jag har funnit nåd för dina ögon, Herre, så må Herren gå med oss. Ty väl är det ett hårdnackat folk, men du vill ju förlåta oss vår missgärning och synd och taga oss till din arvedel.»
Och så skall över eder komma allt rättfärdigt blod som är utgjutet på jorden, ända ifrån den rättfärdige Abels blod intill Sakarias', Barakias' sons blod, hans som I dräpten mellan templet och altaret.
Se, jag skall sända en ängel framför dig, som skall bevara dig på vägen och föra dig till den plats som jag har utsett.
Och det skall ske i kommande dagar att det berg där HERRENS hus är skall stå där fast grundat och vara det yppersta ibland bergen och upphöjt över andra höjder; och alla hednafolk skola strömma dit,
Då stampade hästarnas hovar, när deras tappra ryttare jagade framåt, framåt.
Redan för länge sedan, redan då Saul ännu var konung, var det du som var ledare och anförare för Israel. Och till dig har HERREN, din Gud, sagt: Du skall vara en herde för mitt folk Israel, ja, du skall vara en furste över mitt folk Israel.»
Vi tacka dig, o Gud, vi tacka dig. Ditt namn är oss nära; man förtäljer dina under.
Därefter begav han sig till en stad som hette Nain; och med honom gingo hans lärjungar och mycket folk.
Mose svarade: »Du har talat rätt; jag skall icke vidare komma inför ditt ansikte.»
han som var till i Guds-skepnad, men icke räknade jämlikheten med Gud såsom ett byte,
Men du, människobarn, hör nu vad jag talar till dig; var icke gensträvig såsom detta gensträviga släkte. Öppna din mun och ät vad jag giver dig.»
Och han gav tecken åt dem med handen att de skulle tiga, och förtäljde för dem huru Herren hade fört honom ut ur fängelset. Och han tillade: »Låten Jakob och de andra bröderna få veta detta.» Sedan gick han därifrån och begav sig till en annan ort.
Blevo vi icke av honom aktade såsom främlingar, när han sålde oss? Sedan har han ju ock förtärt vad han fick i betalning för oss.
Sedan vände de båda männen tillbaka och kommo ned från bergsbygden och gingo över floden och kommo så till Josua, Nuns son; och de förtäljde för honom allt vad som hade vederfarits dem.
Och man förde fram sju tjurar, sju vädurar och sju lamm, så ock sju bockar till syndoffer för riket och för helgedomen och för Juda; och han befallde Arons söner, prästerna, att offra detta på HERRENS altare.
Konung Salomo offrade såsom slaktoffer tjugutvå tusen tjurar och ett hundra tjugu tusen av småboskapen. Så invigdes Guds hus av konungen och allt folket.
en uppfostrare för oförståndiga, en lärare för enfaldiga, eftersom du i lagen har uttrycket för kunskapen och sanningen.
Här gäller det för de heliga att hava ståndaktighet, för dem som hålla Guds bud och bevara tron på Jesus.»
Jag skall låta strömmar rinna upp på höjderna och källor i dalarna; jag skall göra öknen till en vattenrik sjö och torrt land till källsprång.
Och i Manasses, Efraims och Simeons städer ända till Naftali genomsökte han överallt husen.
om han ville uppenbara dig sin visdoms lönnligheter, huru han äger förstånd, ja, i dubbelt mått, då insåge du att Gud, dig till förmån, har lämnat åt glömskan en del av din missgärning.
Då sprutade ormen ur sitt gap vatten efter kvinnan såsom en ström, för att strömmen skulle bortföra henne.
Så se nu till; ty HERREN har utvalt dig att bygga ett hus till helgedomen. Var frimodig och gå till verket.»
Och ljusstaken var gjord på följande sätt: den var av guld i drivet arbete; också dess fotställning och blommorna därpå voro i drivet arbete. Efter det mönster som HERREN hade visat Mose hade denne låtit göra ljusstaken.
Men profeten Natan, Benaja, hjältarna och sin broder Salomo inbjöd han icke.
Vidare berättade sekreteraren Safan för konungen och sade: »Prästen Hilkia har givit mig en bok.» Och Safan föreläste den för konungen.
Dessa skaffade sig moabitiska hustrur; den ena hette Orpa och den andra Rut.
vilka hava vågat sina liv för vår Herres, Jesu Kristi, namns skull.
Jag kallade på mina vänner, men de bedrogo mig. Mina präster och mina äldste förgingos i staden, medan de tiggde sig mat för att stilla sin hunger.
Kina, Dimona, Adada,
Och HERREN, din Gud, skall förjaga dessa hedningar för dig, men blott småningom. Du skall icke med hast få förgöra dem, på det att vilddjuren icke må föröka sig till din skada.
gick vidare söder om Skorpionhöjden och fram till Sin, drog sig så upp söder om Kades-Barnea, gick därefter framom Hesron och drog sig upp till Addar samt böjde sig sedan mot Karka.
Och Josef fann nåd för hans ögon och fick betjäna honom. Och han satte honom över sitt hus, och allt vad han ägde lämnade han i hans vård.
Och om han ser ett tåg, ryttare par efter par, ett tåg av åsnor, ett tåg av kameler, då må han giva akt, noga giva akt.»
ty jag säger eder att jag icke mer skall fira denna högtid, förrän den kommer till fullbordan i Guds rike.»
Då svarade han honom: »Välan, jag skall ock häri göra dig till viljes; jag skall icke omstörta den stad som du talar om.
Sådan var den dröm som jag, konung Nebukadnessar, hade. Och du, Beltesassar, må nu säga uttydningen; ty ingen av de vise i mitt rike kan säga mig uttydningen, men du kan det väl, ty heliga gudars ande är i dig.»
Kvinnor funnos som fingo igen sina döda genom deras uppståndelse. Andra läto sig läggas på sträckbänk och ville icke taga emot någon befrielse, i hopp om en så mycket bättre uppståndelse.
Men i konung Joas' tjugutredje regeringsår hade prästerna ännu icke satt i stånd vad som var förfallet på huset.
Och jag skall låta din säd bliva såsom stoftet på jorden; kan någon räkna stoftet på jorden, så skall ock din säd kunna räknas.
Då upptändes Balaks vrede mot Bileam, och han slog ihop händerna. Och Balak sade till Bileam: »Till att förbanna mina fiender kallade jag dig hit, och se, du har i stället nu tre gånger välsignat dem.
och han sover, och han vaknar, och nätter och dagar gå, och säden skjuter upp och växer i höjden, han vet själv icke huru.
Om en man än finge hundra barn och finge leva i många år, ja, om hans livsdagar bleve än så många, men hans själ icke finge njuta sig mätt av hans goda, och om han så bleve utan begravning, då säger jag: lyckligare än han är ett ofullgånget foster.
En livets källa är förståndet för den som äger det, men oförnuftet är de oförnuftigas tuktan.
och färdades genom Syrien och Cilicien och styrkte församlingarna.
Och var och en av eder må taga sitt fyrfat och lägga rökelse därpå, och sedan bära sitt fyrfat fram inför HERRENS ansikte, två hundra femtio fyrfat; du själv och Aron mån ock taga var sitt fyrfat.»
Och David sade till honom: »Ditt blod komme över ditt huvud, ty din egen mun har vittnat mot dig, i det att du sade: 'Jag har dödat HERRENS smorde.'»
Och amoréerna förmådde hålla sig kvar i Har-Heres, Ajalon och Saalbim; men Josefs barns hand blev tung över dem, så att de blevo arbetspliktiga under dessa.
Sen icke därpå att jag är så svart, att solen har bränt mig så. Min moders söner blevo vreda på mig och satte mig till vingårdsvakterska; min egen vingård kunde jag icke vakta.
Böjen edra öron hit och kommen till mig; hören, så får eder själ leva. Jag vill sluta med eder ett evigt förbund: att I skolen undfå all den trofasta nåd jag har lovat David.
Dina präster vare klädda i rättfärdighet, och dina fromma juble.
Och Mose och Aron gjorde alla dessa under inför Farao; men HERREN förstockade Faraos hjärta, så att han icke släppte Israels barn ut ur sitt land.
Och när I kommen in i någon stad där man tager emot eder, så äten vad som sättes fram åt eder,
Förbannen Meros, säger HERRENS ängel, ja, förbannen dess inbyggare, därför att de ej kommo HERREN till hjälp, HERREN till hjälp bland hjältarna.
Så sade nu Gud till Noa: »Detta skall vara tecknet till det förbund som jag har upprättat mellan mig och allt kött på jorden.»
Men när Hiram från Tyrus begav sig ut för att bese de städer som Salomo hade givit honom, behagade de honom icke,
Så säger HERREN: Se, jag skall uppväcka mot Babel och mot Leb-Kamais inbyggare en fördärvares ande.
Därför är jag villig att förkunna evangelium också för eder som bon i Rom.
Och sedan Lemek hade fött Noa, levde han fem hundra nittiofem år och födde söner och döttrar.
Huru förvända ären I icke! Skall då leret aktas lika med krukmakaren? Skall verket säga om sin mästare: »Han har icke gjort mig»? Eller skall bilden säga om honom som har format den: »Han förstår intet»?
Jag skall låta min nitälskan gå över dig, så att de fara grymt fram mot dig; de skola skära av dig näsa och öron, och de som bliva kvar av dig skola falla för svärd. Man skall föra bort dina söner och döttrar, och vad som bliver kvar av dig skall förtäras av eld.
Och somliga läto övertyga sig av det som han sade, men andra trodde icke.
Semaja, Jojarib, Jedaja,
Jag har ofta måst vara ute på resor; jag har utstått faror på floder, faror bland rövare, faror genom landsmän, faror genom hedningar, faror i städer, faror i öknar, faror på havet, faror bland falska bröder --
När sabbaten hade gått till ända, i gryningen till första veckodagen, kommo Maria från Magdala och den andra Maria för att se graven.
Vi hava funnit att denne är en fördärvlig man, som uppväcker strid bland alla judar i hela världen, och att han är en huvudman för nasaréernas parti.
varen såsom jag, som i alla stycken fogar mig efter alla och icke söker min egen nytta, utan de mångas, för att de skola bliva frälsta.
Amrams söner voro Aron och Mose. Och Aron blev jämte sina söner för evärdlig tid avskild till att helgas såsom höghelig, till att för evärdlig tid antända rökelse inför HERREN och göra tjänst inför honom och välsigna i hans namn.
Och framför vaktkamrarna var en avskrankning, som höll en aln; en aln höll ock avskrankningen på motsatta sidan; och var vaktkammare, på vardera sidan, höll sex alnar.
Alltså, mina älskade bröder, varen fasta, orubbliga, alltid överflödande i Herrens verk, eftersom I veten att edert arbete icke är fåfängt i Herren.
och när de nu förnummo vilken nåd som hade blivit mig given, räckte de mig och Barnabas handen till samarbete, både Jakob och Cefas och Johannes, de män som räknades för själva stödjepelarna; vi skulle verka bland hedningarna, och de bland de omskurna.
Och HERREN sade till honom: »Detta är det land som jag med ed har lovat åt Abraham. Isak och Jakob, i det jag sade: 'Åt din säd skall jag giva det.' Jag har nu låtit dig se det med dina ögon, men ditin skall du icke komma.»
När Baal-Hanan, Akbors son, dog, blev Hadar konung efter honom; och hans stad hette Pagu, och hans hustru hette Mehetabel, dotter till Matred, som var dotter till Me-Sahab.
Man bedriver styggelse, var och en med sin nästas hustru; ja, man orenar i skändlighet sin sons hustru; man kränker hos dig sin syster, sin faders dotter.
Och HERRENS ord kom till mig; han sade: Du människobarn, säg till dem:
Strömportarna måste öppna sig, och palatset försmälter av ångest.
utan den plats som HERREN, eder Gud, utväljer inom någon av edra stammar till att där fästa sitt namn, denna boning skolen I söka och dit skall du gå.
Ja, är det icke så med mitt hus inför Gud? Han har ju upprättat med mig ett evigt förbund, i allo stadgat och betryggat. Ja, visst skall han låta all frälsning och glädje växa upp åt mig.
Veten I då icke att de orättfärdiga icke skola få Guds rike till arvedel? Faren icke vilse. Varken otuktiga människor eller avgudadyrkare eller äktenskapsbrytare, varken de som låta bruka sig till synd mot naturen eller de som själva öva sådan synd,
Och han lät leviterna ställa upp sig till tjänstgöring i HERRENS hus med cymbaler, psaltare och harpor, såsom David och Gad, konungens siare, och profeten Natan hade bjudit; ty budet härom var givet av HERREN genom hans profeter.
I de synderna vandraden också I förut, då I ännu haden edert liv i dem.
Konungen frågade honom »Var är han?» Siba svarade konungen: »Han är nu i Makirs, Ammiels sons, hus i Lo-Debar.»
Och härar, utsända av honom, skola komma och oskära helgedomens fäste och avskaffa det dagliga offret och ställa upp förödelsens styggelse.
Här är icke jude eller grek, här är icke träl eller fri, här är icke man och kvinna: alla ären I ett i Kristus Jesus.
Kraftverkningarna äro mångahanda, men Gud är en och densamme, han som verkar allt i alla.
Lyft det sedan i deras åsyn upp på axeln och för bort det, när det har blivit alldeles mörkt; och betäck ditt ansikte, så att du icke ser landet. Ty jag gör dig till ett tecken för Israels hus.»
Då sade jag till min herre: 'Men om nu kvinnan icke vill följa med mig?'
allt såsom HERREN hade bjudit Mose; och han mönstrade dem i Sinais öken.
Hans huvud och hår var vitt såsom vit ull, såsom snö, och hans ögon voro såsom eldslågor.
Men männen ville icke höra på honom; då tog mannen sin bihustru och förde henne ut till dem. Och de kände henne och hanterade henne skändligt hela natten ända till morgonen; först när morgonrodnaden gick upp, läto de henne gå.
»Dessa voro de män från hövdingdömet, som drogo upp ur den landsflykt och fångenskap till vilken de hade blivit bortförda av Nebukadnessar, konungen i Babel, och som vände tillbaka till Jerusalem och till Juda, var och en till sin stad,
Huru skall en yngling bevara sin väg obesmittad? När han håller sig efter ditt ord.
Den som har öra, han höre vad Anden säger till församlingarna.»
Och Faraos dotter kom ned till floden för att bada, och hennes tärnor gingo utmed floden. När hon nu fick se kistan i vassen, sände hon sin tjänarinna dit och lät hämta den till sig.
Alla dessa höllo endräktigt ut i bön tillika med Maria, Jesu moder, och några andra kvinnor samt Jesu bröder.
Och Saul och allt det folk som han hade hos sig församlade sig och drogo till stridsplatsen; där fingo de se att den ene hade lyft sitt svärd mot den andre, så att en mycket stor förvirring hade uppstått.
Ty jag är viss om att varken död eller liv, varken änglar eller andefurstar, varken något som nu är eller något som skall komma,
Det må vara lärjungen nog, om det går honom såsom hans mästare, och tjänaren, om det går honom såsom hans herre. Om de hava kallat husbonden för Beelsebul, huru mycket mer skola de icke så kalla hans husfolk!
Därför säger HERREN så om Anatots män, dem som stå efter ditt liv och säga: »Profetera icke i HERRENS namn, om du icke vill dö för vår hand»
Sedan trädde de fram till honom och sade: »Hell dig, du judarnas konung!» och slogo honom på kinden.
åt denne inrett en stor kammare, där man förut plägade lägga in spisoffret, rökelsen och kärlen och den tionde av säd, vin och olja, som var bestämd åt leviterna, sångarna och dörrvaktarna, så ock offergärden åt prästerna.
Ja, alla andra folk vandra vart och ett i sin guds namn, men vi vilja vandra i HERRENS, vår Guds, namn, alltid och evinnerligen.
När lärjungarna sågo detta, förundrade de sig och sade: »Huru kunde fikonträdet så i hast förtorkas?»
Och prästerna, Levi söner, skola träda fram, ty dem har HERREN, din Gud, utvalt till att göra tjänst inför honom och till att välsigna i HERRENS namn, och såsom de bestämma skola alla tvister och alla misshandlingsmål behandlas.
Så ofta israeliterna hade sått, drogo midjaniterna, amalekiterna och österlänningarna upp emot dem
Vid deras åsyn gripas folken av ångest, alla ansikten skifta färg.
Och Aron var ett hundra tjugutre år gammal, när han dog på berget Hor.
I samma stund kommo några fariséer fram och sade till honom: »Begiv dig åstad bort härifrån; ty Herodes vill dräpa dig.»
Och han förde fram brännoffersväduren, och Aron och hans söner lade sina händer på vädurens huvud.
Då trädde en av de skriftlärde fram, en som hade hört deras ordskifte och förstått att han hade svarat dem väl. Denne frågade honom: »Vilket är det förnämsta av alla buden?»
Eftersom I genom lögnaktigt tal haven gjort den rättfärdige försagd i hjärtat, honom som jag ingalunda ville plåga, men däremot haven styrkt den ogudaktiges mod, så att han icke vänder om från sin onda väg och räddar sitt liv,
Men alltsammans kommer från Gud, som har försonat oss med sig själv genom Kristus och givit åt oss försoningens ämbete.
Men jag hämtade eder fader Abraham från andra sidan floden och lät honom vandra omkring i hela Kanaans land. Och jag gjorde hans säd talrik; jag gav honom Isak,
Och Farao blev förtörnad på sina två hovmän, överste munskänken och överste bagaren,
Då nu Jesus märkte att han hade svarat förståndigt, sade han till honom: »Du är icke långt ifrån Guds rike.» Sedan dristade sig ingen att vidare ställa någon fråga på honom.
och sade: »Herre, min tjänare ligger därhemma lam och lider svårt.»
Då svarade allt folket med en mun och sade: »Allt vad HERREN har talat vilja vi göra.» Och Mose gick tillbaka till HERREN med folkets svar.
Och om ditt offer är ett spisoffer som tillredes på plåt, så skall det vara av fint mjöl, begjutet med olja, osyrat.
och de talade inställsamt för honom med sin mun och skrymtade för honom med sin tunga.
Om han vill bära fram ett brännoffer av fäkreaturen, så skall han därtill taga ett felfritt djur av hankön och föra det fram till uppenbarelsetältets ingång, för att han må bliva välbehaglig inför HERRENS ansikte.
På samma sätt hade han gjort för Esaus barn, som bo i Seir, i det han för dem förgjorde horéerna; de fördrevo dem och bosatte sig i deras land, där de bo ännu i dag.
Det bud som Jonadab, Rekabs son, gav sina barn, att de icke skulle dricka vin, det har blivit iakttaget, och ännu i dag dricka de icke vin, av hörsamhet mot sin faders bud. Men själv har jag titt och ofta talat till eder, och I haven dock icke hörsammat mig.
Och däri består kärleken, att vi vandra efter de bud han har givit. Ja, detta är budet, att I skolen vandra i kärleken, enligt vad I haven hört från begynnelsen.
Hon bliver ock agad genom plågor på sitt läger och genom ständig oro, allt intill benen.
Gören därför bättring och omvänden eder, så att edra synder bliva utplånade,
Men där var ock en annan stor örn med stora vingar och fjädrar i mängd; och se, till denne böjde nu vinträdet längtansfullt sina grenar, och från platsen där det var planterat sträckte det sina rankor mot honom, för att han skulle vattna det.
Jag vill höra vad Gud, HERREN, talar: se, han talar frid till sitt folk och till sina fromma; må de blott icke vända åter till dårskap.
Och hövding för gersoniternas stamfamilj var Eljasaf, Laels son.
Ty då hedningarna, som icke hava lag, av naturen göra vad lagen innehåller, så äro dessa, utan att hava lag, sig själv en lag,
Och konung David sade till hela församlingen: »Min son Salomo den ende som Gud har utvalt, är ung och späd, och arbetet är stort, ty denna borg är icke avsedd för en människa, utan för HERREN Gud.
Då nu Jesus märkte att han hade svarat förståndigt, sade han till honom: »Du är icke långt ifrån Guds rike.» Sedan dristade sig ingen att vidare ställa någon fråga på honom.
Och Mose och Aron och hans söner tvådde sedermera sina händer och fötter med vatten därur;
»Sannerligen, sannerligen säger jag eder: Den som icke går in i fårahuset genom dörren, utan stiger in någon annan väg, han är en tjuv och en rövare.
Den som ävlas att få vänner, han kommer i olycka; men vänner finnas, mer trogna än en broder.
hans offergåva var ett silverfat, ett hundra trettio siklar i vikt, och en silverskål om sjuttio siklar, efter helgedomssikelns vikt, båda fulla med fint mjöl, begjutet med olja, till spisoffer,
Genom att höra på dem förökar den vise sin lärdom och förvärvar den förståndige rådklokhet.
Och du, människobarn, profetera Och såg: Så säger Herren, HERREN om Ammons barn och om deras smädelser: Säg: Ett svärd, ja, ett svärd är draget, det är fejat för att slakta för att varda mättat och för att blixtra,
Därför skall deras väg bliva för dem såsom en slipprig stig i mörkret, de skola på den stöta emot och falla. Ty jag vill låta olycka drabba dem, när deras hemsökelses är kommer, säger HERREN.
Låten båda slagen växa tillsammans intill skördetiden; och när skördetiden är inne, vill jag säga till skördemännen: 'Samlen först tillhopa ogräset, och binden det i knippor till att brännas upp, och samlen sedan in vetet i min lada.'»
Men de ropade till HERREN i sin nöd, och han frälste dem ur deras trångmål;
Det lilla som en rättfärdig har är bättre än många ogudaktigas stora håvor.
Det är icke I som skolen tala, utan det är eder Faders Ande som skall tala i eder.
Och HERREN bjöd oss att göra efter all dessa stadgar och att frukta HERREN, vår Gud, för att det alltid skulle gå oss väl, i det att han behölle oss vid liv, såsom ock hittills har skett.
Och Gud välsignade dem; Gud sade till dem: »Varen fruktsamma och föröken eder, och uppfyllen jorden och läggen den under eder; och råden över fiskarna i havet och över fåglarna under himmelen och över alla djur som röra sig på jorden.»
Dina heliga städer hava blivit en öken, Sion har blivit en öken, Jerusalem en ödemark.
Och han lät oss komma hit och gav oss detta land, ett land som flyter av mjölk och honung.
Om nu Satan driver ut Satan, så har han kommit i strid med sig själv. Huru kan då hans rike hava bestånd?
Så föllo av Benjamin aderton tusen man, allasammans tappert folk.
Och vad du måste utbetala för det som härutöver behöves till din Guds hus, det må du låta utbetala ur konungens skattkammare.
Tjänen HERREN med glädje, kommen inför hans ansikte med fröjderop.
Och ur korgen med de osyrade bröden, som stod inför HERRENS ansikte, tog han en osyrad kaka, en oljebrödskaka och en tunnkaka och lade detta på fettstyckena och det högra lårstycket.
Och fönster funnos på den och på dess förhus runt omkring, likadana som de andra fönstren. Den var femtio alnar lång och tjugufem alnar bred.
Ja, klagoropen ljuda runtom i Moabs land; till Eglaim når dess jämmer och till Beer-Elim dess jämmer.
utan du skall gå till den plats som Herren, din Gud, utväljer till boning åt sitt namn, och där skall du slakta påskoffret om aftonen, när solen går ned den tid på dagen, då den drog ut ur Egypten.
Ty en annan grund kan ingen lägga, än den som är lagd, nämligen Jesus Kristus;
Och ingen annan rökelse mån I göra åt eder så sammansatt som denna skall vara. Helig skall den vara dig för HERREN.
Och striden blev på den dagen allt häftigare, och Israels konung höll sig ända till aftonen upprätt i sin vagn, vänd mot araméerna; men vid den tid då solen gick ned gav han upp andan.
Vaken, och bedjen att I icke mån komma i frestelse. Anden är villig, men köttet är svagt.»
Då svarade Jesus honom: »Rävarna hava kulor, och himmelens fåglar hava nästen; men Människosonen har ingen plats där han kan vila sitt huvud.»
Ett falskt vittne bliver icke ostraffat, och den som främjar lögn, han kommer icke undan.
Likväl sänder jag nu åstad dessa bröder, för att det som jag har sagt till eder berömmelse icke skall i denna del befinnas hava varit tomt tal. Ty, såsom jag förut har sagt, jag vill att I skolen vara redo.
Kallar jag på min tjänare, så svarar han icke; ödmjukt måste jag bönfalla hos honom.
Och över judarnas äldste vakade deras Guds öga, så att man lovade att icke lägga något hinder i vägen för dem, till dess saken hade kommit inför Darejaves; sedan skulle man sända dem en skrivelse härom.
Konungen frågade: »Finnes ingen kvar av Sauls hus, mot vilken jag kan bevisa barmhärtighet, såsom Gud är barmhärtig?» Siba svarade konungen: »Ännu finnes kvar en son till Jonatan, en som är ofärdig i fötterna.»
han höll nämligen Kristi smälek för en större rikedom än Egyptens skatter, ty han hade sin blick riktad på lönen.
ty du vet att en sådan är förvänd och begår synd, ja, han har själv fällt domen över sig.
Den som fruktar HERREN, han vandrar i redlighet, men den som föraktar honom, han går krokiga vägar.
Väduren som du såg, han med de två hornen, betyder Mediens och Persiens konungar.
Där uppehöll han sig i tre månader. När han sedan tänkte avsegla därifrån till Syrien, beslöt han, eftersom judarna förehade något anslag mot honom, att göra återfärden genom Macedonien.
Och överhovmästaren Eljakim och sekreteraren Sebna och de äldste bland prästerna sände han, höljda i sorgdräkt, till profeten Jesaja, Amos' son.
Och du skall göra femtio häktor av guld och foga tillhopa våderna med varandra medelst häktorna, så att tabernaklet utgör ett helt.
och sade: »Så skolen I säga: 'Hans lärjungar kommo om natten och stulo bort honom, medan vi sovo.'
Av den minste skola komma tusen, och av den ringaste skall bliva ett talrikt folk. Jag är HERREN; när tiden är inne, skall jag med hast fullborda detta.
Och de bådo och sade: »Herre, du som känner allas hjärtan, visa oss vilken av dessa två du har utvalt
bjöd han leviterna som buro HERRENS förbundsark och sade:
Gören därför bättring och omvänden eder, så att edra synder bliva utplånade,
Ty väl är det fåfängt, då man vill fånga fåglar, att breda ut nätet i hela flockens åsyn.
Och var och en som icke gör efter din Guds lag och konungens lag, över honom skall dom fällas med rättvisa, vare sig till död eller till landsförvisning eller till penningböter eller till fängelse.»
Ja, förstår du himmelens lagar, och ordnar du dess välde över jorden?
Men de stodo stilla, var och en på sin plats, runt omkring lägret. Då begynte alla i lägret att löpa hit och dit och skria och fly.
Må deras bord framför dem bliva till en snara och till ett giller, bäst de gå där säkra;
Det har blivit ditt fördärv, o Israel, att du satte dig upp mot mig som var din hjälp.
Men Jonatan, Davids farbroder, var rådgivare; han var en förståndig och skriftlärd man. Jehiel, Hakmonis son, var anställd hos konungens söner.
av Josefs barn: av Efraim: Elisama, Ammihuds son; av Manasse: Gamliel, Pedasurs son;
fick han fatt på en ung man, en av invånarna i Suckot, och utfrågade denne, och han måste skriva upp åt honom de överste i Suckot och de äldste där, sjuttiosju män.
Och Hosea, Elas son, anstiftade en sammansvärjning mot Peka, Remaljas son, och slog honom till döds och blev så konung i hans ställe, i Jotams, Ussias sons, tjugonde regeringsår.
Men kaldéernas här förföljde konungen, och de hunno upp honom på Jerikos hedmarker, sedan hela hans här hade övergivit honom och skingrat sig.
Ty var och en som beder, han får; och den som söker, han finner; och för den som klappar skall varda upplåtet.
Du skall trolova dig med en kvinna, men en annan man skall sova hos henne; du skall bygga ett hus, men icke få bo däri; du skall plantera en vingård, men icke få skörda dess frukt.
Om jag nu har anbefallt Titus, så mån I besinna att han är min medbroder och min medarbetare till edert bästa; och om jag har skrivit om andra våra bröder, så mån I besinna att de äro församlingssändebud och Kristi ära.
Eftersom du är så dyrbar i mina ögon, så högt aktad och så älskad av mig, därför giver jag människor till lösen för dig och folk till lösen för ditt liv.
Mina sabbater skolen I hålla, och för min helgedom skolen I hava fruktan. Jag är HERREN.
hedningarna åter hava fått prisa Gud för hans barmhärtighets skull. Så är ock skrivet: »Fördenskull vill jag prisa dig bland hedningarna och lovsjunga ditt namn.»
Ditt majestäts härlighet och ära vill jag begrunda och dina underfulla verk.
Men somt föll i god jord, och det sköt upp och växte och gav frukt och bar trettiofalt och sextiofalt och hundrafalt.»
Men när han hörde detta, blev han djupt bedrövad, ty han var mycket rik.
Vad orsak haven I till att bruka detta ordspråk i Israels land: »Fäderna äta sura druvor, och barnens tänder bliva ömma därav»?
Och Jakob flydde till Arams mark Israel tjänade för en kvinna, för en kvinnas skull vaktade han hjorden.
Och han kom tillbaka till Juda och sade: »Jag har icke funnit henne; därtill säger folket på orten att ingen tempeltärna har varit där.»
Det har varit för mig en stor glädje i Herren att I nu omsider haven kommit i en så god ställning, att I haven kunnat tänka på mitt bästa. Dock, I tänkten nog också förut därpå, men I haden icke tillfälle att göra något.
Kus' söner voro Seba, Havila, Sabta, Raema och Sabteka. Raemas söner voro Saba och Dedan.
Uppe på höjderna står hon, vid vägen, där stigarna mötas.
Om någon icke vill omvända sig, så vässer han sitt svärd, sin båge spänner han och gör den redo;
Esau sade till sin fader: »Har du då allenast den enda välsignelsen, min fader? Välsigna också mig, min fader.» Och Esau brast ut i gråt.
HERREN är sitt folks starkhet, och ett frälsningens värn är han för sin smorde.
Då han emellertid ville få säkert besked om varför Paulus anklagades av judarna, låt han dagen därefter taga av honom bojorna och bjöd översteprästerna och hela Stora rådet att komma tillsammans. Sedan lät han föra Paulus ditned och ställde honom inför dem.
Om en prästs dotter ohelgar sig genom skökolevnad, så ohelgar hon sin fader; hon skall brännas upp i eld.
fattade hon honom i manteln och sade: »Ligg hos mig.» Men han lämnade manteln i hennes hand och flydde och kom ut.
Då sade han till honom: »Eftersom du icke har lyssnat till HERRENS röst, därför skall ett lejon slå ned dig, när du går ifrån mig.» Och när han gick sin väg ifrån honom, kom ett lejon emot honom och slog ned honom.
ej heller skall du i ditt hus hava två slags efa-mått, ett större och ett mindre.
Folket, som stod där och hörde detta, sade då: »Det var ett tordön.» Andra sade: »Det var en ängel som talade med honom.»
Sion hör det och gläder sig, och Juda döttrar fröjda sig för dina domars skull, HERRE.
Här visade sig för Paulus i en syn om natten en macedonisk man, som stod där och bad honom och sade: »Far över till Macedonien och hjälp oss.»
Upp, alla I som ären törstiga, kommen hit och fån vatten; och I som inga penningar haven, kommen hit och hämten säd och äten. Ja, kommen hit och hämten säd utan penningar och för intet både vin och mjölk.
Tänk, min Gud på Tobia, ävensom Sanballat, efter dessa hans gärningar, så ock på profetissan Noadja och de andra profeterna som ville skrämma mig!
Men jag har något litet emot dig: du har hos dig några som hålla fast vid Balaams lära, hans som lärde Balak huru han skulle lägga en stötesten för Israels barn, så att de skulle äta kött från avgudaoffer och bedriva otukt.
Då nu Moses svärfader såg allt vad han hade att beställa med folket, sade han: »Vad är det allt du har att bestyra med folket? Varför sitter du här till doms ensam under det att allt folket måste stå omkring dig från morgonen ända till aftonen?»
För sångmästaren; av Koras söner; en psalm.
Ty deras vredes stora dag är kommen, och vem kan bestå?»
Och Hiskia gick till vila hos sina fäder. Och hans son Manasse blev konung efter honom.
Och till Amasa skolen I säga: 'Är du icke mitt kött och ben? Gud straffe mig nu och framgent, om du icke för all din tid skall bliva härhövitsman hos mig i Joabs ställe.'»
Så skall då Herren, HERREN Sebaot sända tärande sjukdom i hans feta kropp, och under hans härlighet skall brinna en brand likasom en brinnande eld.
Ty dessa lade alla dit av sitt överflöd, men hon lade dit av sitt armod allt vad hon hade, så mycket som fanns i hennes ägo.»
Och de fem män som hade varit åstad för att bespeja landet gingo upp och kommo ditin och togo den skurna gudabilden och efoden, så ock husgudarna och den gjutna gudabilden, under det att prästen stod vid ingången till porten jämte de sex hundra vapenomgjordade männen.
Jag levde en gång utan lag; men när budordet kom, fick synden liv,
Vi älska dem för sanningens skull, som förbliver i oss, och som skall vara med oss till evig tid.
Detta är vad som stod i det brev som profeten Jeremia sände från Jerusalem till de äldste som ännu levde kvar i fångenskapen, och till prästerna och profeterna och allt folket, dem som Nebukadnessar hade fört bort ifrån Jerusalem till Babel,
Förhuset var tjugu alnar lång och elva alnar brett, nämligen vid trappstegen på vilka man steg ditupp. Och vid murpelarna stodo pelare, en på var sida.
När Hirams flotta hämtade guld från Ofir, hemförde också den från Ofir almugträ i stor myckenhet, ävensom ädla stenar.
Skära mig med isop, så att jag varder ren; två mig, så att jag bliver vitare än snö.
Ty det ordet skulle fullbordas, som han hade sagt: »Av dem som du har givit mig har jag icke förlorat någon.»
239400
En bihustru som han hade i Sikem födde honom ock en son; denne gav han namnet Abimelek.
Icke är jag väl ett hav eller ett havsvidunder, så att du måste sätta ut vakt mot mig?
Låt varna dig, Jerusalem, så att min själ ej vänder sig ifrån dig, så att jag icke gör dig till en ödemark, till ett obebott land.
Och Jesus talade till honom och sade: »Vad vill du att jag skall göra dig?» Den blinde svarade honom: »Rabbuni, låt mig få min syn.»
Ben-Geber i Ramot i Gilead; han hade Manasses son Jairs byar, som ligga i Gilead; han hade ock landsträckan Argob, som ligger i Basan, sextio stora städer med murar och kopparbommar;
Och du skall älska HERREN, din Gud, av allt ditt hjärta och av all din själ och av all din kraft.
Och Jakob sade till sina fränder: »Samlen tillhopa stenar.» Och de togo stenar och gjorde ett röse och höllo måltid där på röset.
Om däremot någon är fast i sitt sinne och icke bindes av något nödtvång, utan kan följa sin egen vilja, och så i sitt sinne är besluten att låta sin ogifta dotter förbliva såsom hon är, då gör denne väl.
Och den som skall renas skall två sina kläder och raka av allt sitt hår och bada sig i vatten, så bliver han ren och får sedan gå in i lägret. Dock skall han stanna utanför sitt tält i sju dagar.
De svulster av guld som filistéerna gåvo såsom skuldoffer åt HERREN utgjorde: för Asdod en, för Gasa en, för Askelon en, för Gat en, för Ekron en.
Och Johannes hade kläder av kamelhår och bar en lädergördel om sina länder och levde av gräshoppor och vildhonung.
Ställ dig i porten till HERRENS hus, och predika där detta ord och säg: Hören HERRENS ord, I alla av Juda, som gån in genom dessa portar för att tillbedja HERREN.
När Saul nu hade tagit konungadömet över Israel i besittning, förde han krig mot alla sina fiender runt omkring: mot Moab, mot Ammons barn, mot Edom, mot konungarna i Soba och mot filistéerna; och vart han vände sig tuktade han dem.
Och Josef dog, när han var ett hundra tio år gammal. Och man balsamerade honom, och han lades i en kista, i Egypten.
aviterna gjorde sig en Nibhas och en Tartak, och sefarviterna brände upp sina barn i eld åt Adrammelek och Anammelek, Sefarvaims gudar.
De befästa sig i sitt onda uppsåt, de orda om huru de skola lägga ut snaror; de säga: »Vem skulle se oss?»
varhelst någon oförvitlig man funnes, en enda kvinnas man, en som hade troende barn, vilka icke vore i vanrykte för oskickligt leverne eller vore uppstudsiga.
Och den omfattade Kattat, Nahalal, Simron, Jidala och Bet-Lehem -- tolv städer med deras byar.
Mjölk gav jag eder att dricka; fast föda gav jag eder icke, ty det fördrogen I då ännu icke. Ja, icke ens nu fördragen I det,
Därför säger Herren, HERREN så: Eftersom edert tal är falskhet och edra syner äro lögn, se, därför skall jag komma över eder, säger Herren, HERREN.
Och HERRENS tjänare Mose dog där i Moabs land, såsom HERREN hade sagt.
Ty ljusets frukt består i allt vad godhet och rättfärdighet och sanning är.
Och när folket såg honom, lovade de likaledes sin gud och sade: »Vår gud har givit vår fiende i vår hand honom som förödde vårt land och slog så många av oss ihjäl.»
När de hörde detta, prisade de Gud. Och de sade till honom: »Du ser, käre broder, huru många tusen judar det är som hava kommit till tro, och alla nitälska de för lagen.
Lottkastning gör en ände på trätor, den skiljer mellan mäktiga män.
Visserligen har allt detta fått namn om sig att vara »vishet», eftersom däri ligger ett självvalt gudstjänstväsende och ett slags »ödmjukhet» och en kroppens späkning; men ingalunda ligger däri »en viss heder», det tjänar allenast till att nära det köttsliga sinnet.
Då svarade Jakob och sade till Laban: »Jag fruktade för dig, ty jag tänkte att du skulle med våld taga dina döttrar ifrån mig.
Då drog konung Joram ut från Samaria och mönstrade hela Israel.
HERREN är konung evinnerligen, din Gud, Sion, från släkte till släkte. Halleluja!
Men staden med allt vad däri är skall givas till spillo åt HERREN; allenast skökan Rahab skall få leva, jämte alla som äro inne i hennes hus, därför att hon gömde de utskickade som vi hade sänt åstad.
så många av Efraims stam som inmönstrades; utgjorde fyrtio tusen fem hundra.
Men över Davids hus och över Jerusalems invånare skall jag utgjuta en nådens och bönens ande, så att de se upp till mig, och se vem de hava stungit. Och de skola hålla dödsklagan efter honom, såsom man håller dödsklagan efter ende sonen, och skola bittert sörja honom, såsom man sörjer sin förstfödde.
Åter talade Jesus till dem och sade: »Jag är världens ljus; den som följer mig, han skall förvisso icke vandra i mörkret, utan skall hava livets ljus.»
Tagen därför ifrån honom hans pund, och given det åt den som har de tio punden.
Eller är Gud allenast judarnas Gud? Är han icke ock hedningarnas? Jo, förvisso också hedningarnas,
I världen var han, och genom honom hade världen blivit till, men världen ville icke veta av honom.
Så låtom oss lära känna HERREN, ja, låtom oss fara efter att lära känna honom. Hans uppgång är så viss som morgonrodnadens, och han skall komma över oss lik ett regn, lik ett vårregn, som vattnar jorden.»
Åt denne gav då Simon Petrus ett tecken och sade till honom: »Säg vilken det är som han talar om.»
så många av Naftali stam som inmönstrades, utgjorde femtiotre tusen fyra hundra.
Rök steg upp från hans näsa och förtärande eld från hans mun; eldsglöd ljungade från honom.
Inom sina förtryckares murar måste de bereda olja, de få trampa vinpressar och därvid lida törst.
Och Abram blev av honom väl behandlad för hennes skull, så att han fick får, fäkreatur och åsnor, tjänare och tjänarinnor, åsninnor och kameler.
Gåvor öppna väg för en människa och föra henne fram inför de store.
Nej, I gören eder faders gärningar.» De sade till honom: »Vi äro icke födda i äktenskapsbrott. Vi hava Gud till fader och ingen annan.»
Och jag skall sätta dem till att förrätta tjänsten i huset vid allt tjänararbete där, allt som där skall utföras.
Därför, om nu en profet profeterar om lycka, så kan man först då när den profetens ord går i fullbordan veta att han är en profet som HERREN i sanning har sänt.»
Och edra altaren skola varda förödda och edra solstoder sönderkrossade, och dem av eder, som bliva slagna, skall jag låta bliva kastade inför edra eländiga avgudar.
Mosa födde Binea. Hans son var Rafa; hans son var Eleasa; hans son var Asel.
Om någon ligger hos sin svärdotter, så skola de båda straffas med döden; de hava bedrivit en vederstygglighet, blodskuld låder vid dem.
Jag sade i mitt hjärta: »Se, jag har förvärvat mig stor vishet, och jag har förökat den, så att den övergår allas som före mig hava regerat över Jerusalem; ja, vishet och insikt har mitt hjärta inhämtat i rikt mått.»
Men när Cefas kom till Antiokia, trädde jag öppet upp mot honom, ty han hade befunnits skyldig till en försyndelse.
då skall du överlämna åt HERREN allt det som öppnar moderlivet. Allt som öppnar moderlivet av det som födes bland din boskap skall, om det är hankön, höra HERREN till.
så att markens djur skola ära mig, schakaler och strutsar, därför att jag låter vatten flyta i öknen, strömmar i ödemarken, så att mitt folk, min utkorade, kan få dricka.
Där fanns nämligen en guldsmed, vid namn Demetrius, som förfärdigade Dianatempel av silver och därmed skaffade hantverkarna en ganska stor inkomst.
Skapa i mig, Gud, ett rent hjärta, och giv mig på nytt en frimodig ande.
Och ännu mycket tydligare blir detta, då nu en präst av annat slag uppstår, lik Melkisedek däri,
Ty alla de som drivas av Guds Ande, de äro Guds barn.
David själv har ju sagt genom den helige Andes ingivelse: 'Herren sade till min herre: Sätt dig på min högra sida, till dess jag har lagt dina fiender dig till en fotapall.'
Om du framlägger detta för bröderna, så bevisar du dig såsom en god Kristi Jesu tjänare, då du ju hämtar din näring av trons och den goda lärans ord, den läras som du troget har efterföljt.
och vinnläggen eder om att bevara Andens enhet genom fridens band:
Därifrån gick den fram österut mot solens uppgång till Gat-Hefer och Et-Kasin och vidare till det Rimmon som sträcker sig till Nea.
då när Gud stod upp till dom, till att frälsa alla ödmjuka på jorden. Sela.
och i vilken man såg profeters och heliga mäns blod, ja, alla de människors blod, som hade blivit slaktade på jorden.»
När han sedan lät Benjamins stam gå fram efter dess släkter, träffade Matris släkt av lotten; därpå träffades Saul, Kis' son, av lotten, men när de då sökte efter honom, stod han icke att finna.
I veten ju vilka bud vi hava givit eder genom Herren Jesus.
Vem mäktar rycka av honom hans pansar? Vem vågar sig in mellan hans käkars par?
Där må prästen Sadok och profeten Natan smörja honom till konung över Israel; sedan skolen I stöta i basun och ropa: 'Leve konung Salomo!'
Och somt föll på stengrund, och när det hade vuxit upp, torkade det bort, eftersom det icke där hade någon fuktighet.
Du gör oss till ett trätoämne för våra grannar, och våra fiender bespotta oss.
Nåd vare med eder och frid ifrån Gud, Fadern, och Herren Jesus Kristus.
Jag skall bliva för Israel såsom dagg, han skall blomstra såsom en lilja, och såsom Libanons skog skall han skjuta rötter.
Därför säger HERREN så om konungen i Assyrien: Han skall icke komma in i denna stad och icke skjuta någon pil ditin; han skall icke mot den föra fram någon sköld eller kasta upp någon vall mot den.
Giv mig, min son, ditt hjärta, och låt mina vägar behaga dina ögon.
Bileam, Beors son, spåmannen, dräptes ock av Israels barn med svärd, jämte andra som då blevo slagna av dem.
Därför säger Herren, HERREN Sebaot så: Frukta icke, mitt folk, du som bor i Sion, för Assur, när han slår dig med riset och upplyfter sin stav mot dig, såsom man gjorde i Egypten.
När då Husai kom in till Absalom, sade Absalom till honom: »Så och så har Ahitofel talat. »Skola vi göra såsom han har sagt? Varom icke, så tala du.»
Hör, dottern mitt folk ropar i fjärran land: »Finnes då icke HERREN i Sion? Är dennes konung icke mer där?» Ja, varför hava de förtörnat mig med sina beläten, med sina främmande avgudar?
Och i din vingård skall du icke göra någon efterskörd, och de avfallna druvorna i din vingård skall du icke plocka upp; du skall lämna detta kvar åt den fattige och åt främlingen. Jag är HERREN, eder Gud.
Att man krossar under sina fötter alla fångar i landet,
I åter skolen icke sluta förbund med detta lands inbyggare; I skolen bryta ned deras altaren.' Men I haven icke velat höra min röst. Vad haven I gjort! --
den femtonde lotten kom ut för Jeremot, med hans söner och bröder, tillsammans tolv;
och talen till varandra i psalmer och lovsånger och andliga visor, och sjungen och spelen till Herrens ära i edra hjärtan,
Och när Jehu kom in genom porten, ropade hon: »Allt står väl rätt till, du, Simri, som har dräpt din herre?»
Och HERREN har i dag hört dig förklara att du vill vara hans egendomsfolk, såsom han har sagt till dig, och att du vill hålla alla hans bud;
Sedan begav han sig åstad till Tarsus för att uppsöka Saulus.
Och Samuel tog sin oljeflaska och göt olja på hans huvud och kysste honom och sade: »Se, HERREN har smort dig till furste över sin arvedel.
Och Darejaves av Medien mottog riket, när han var sextiotvå år gammal.
Hans ben äro pelare av vitaste marmor, som vila på fotstycken av finaste guld. Att se honom är såsom att se Libanon; ståtlig är han såsom en ceder.
Ty deras bördeman är stark; han skall utföra deras sak mot dig.
Och prästerna, leviterna, dörrvaktarna, sångarna, en del av meniga folket samt tempelträlarna, korteligen hela Israel, bosatte sig i sina städer.»
Herren låter höra sitt ord, stor är skaran av kvinnor som båda glädje:
Och Josef sade till sina bröder: »Jag dör, men Gud skall förvisso se till eder, och föra eder upp från detta land till det land som han med ed har lovat åt Abraham, Isak och Jakob.»
Rikligen mättad är vår själ med de säkras bespottelse, med de högmodigas förakt.
Denna sade till sin fru: »Ack att min herre vore hos profeten i Samaria, så skulle denne nog befria honom från hans spetälska!»
så kan det grönska upp genom vattnets ångor och skjuta grenar lik ett nyplantat träd.
Åtta dagar därefter voro hans lärjungar åter därinne, och Tomas var med bland dem. Då kom Jesus, medan dörrarna voro stängda, och stod mitt ibland de, och sade: »Frid vare med eder!»
då skall du svara din son: »Vi voro Faraos trälar i Egypten, men med stark hand förde HERREN oss ut ur Egypten.
Men en tjänstekvinna, som fick se honom, där han satt vid elden fäste ögonen på honom och sade: »Också denne var med honom.
Och en man i folkhopen svarade honom: »Mästare, jag har fört till dig min son, som är besatt av en stum ande.
Men om en ängel då finnes, som vakar över henne, en medlare, någon enda av de tusen, och denne får lära människan hennes plikt,
Vad man nu därutöver söker hos förvaltare är att en sådan må befinnas vara trogen.
Min insikt vill jag hämta vida ifrån, och åt min skapare vill jag skaffa rätt.
Voren I av världen, så älskade ju världen vad henne tillhörde; men eftersom I icke ären av världen, utan av mig haven blivit utvalda och tagna ut ur världen, därför hatar världen eder.
säg: Hör HERRENS ord, du Juda konung, som sitter på Davids tron, hör det du med dina tjänare och ditt folk, I som gån in genom dessa portar.
Och han kom till den andre och sade sammalunda. Då svarade denne och sade: 'Ja, herre'; men han gick icke,
Då sade hon: »Se, din svägerska har vänt tillbaka till sitt folk och till sin gud; vänd ock du tillbaka och följ din svägerska.»
Och allt folket och hela Israel insåg då att konungen ingen del hade haft i att Abner, Ners son, hade blivit dödad.
Och Jesus sade: »Till en dom har jag kommit hit i världen, för att de som icke se skola varda seende, och för att de som se skola varda blinda.»
Och detta är lagen om skuldoffret: Det är högheligt.
Och jag skall föra Israel tillbaka till hans betesmarker, och han skall få gå bet på Karmel och i Basan; och på Efraims berg och i Gilead skall han få äta sig mätt.
Sjungen till hans ära, lovsägen honom, talen om alla hans under.
eller i det att han, när han har hittat något borttappat, nekar därtill och svär falskt i någon sak, vad det nu må vara, vari en människa kan försynda sig:
Av en talent rent guld skall man göra den med alla dessa tillbehör.
De skola sjunga om HERRENS vägar, ty HERRENS ära är stor.
med nardus och saffran, kalmus och kanel och rökelseträd av alla slag, med myrra och aloe och de yppersta kryddor av alla slag.
När bröderna förnummo detta, förde de honom ned till Cesarea och sände honom därifrån vidare till Tarsus.
Foga dem sedan tillhopa med varandra till en enda stav, så att de bliva förenade till ett i din hand.
Jesus svarade och sade till dem: »Om jag än vittnar om mig själv, så gäller dock mitt vittnesbörd, ty jag vet varifrån jag har kommit, och vart jag går; men I veten icke varifrån jag kommer, eller vart jag går.
Käre bröder, bedjen för oss.
Men lika lätt kan en dåraktig man få förstånd, som en vildåsnefåle kan födas till människa.
Huru länge, HERRE, skall jag ropa, utan att du hör klaga inför dig över våld, utan att du frälsar?
Då sade han till dem: »Från storätaren utgick ätbart, från den grymme kom sötma.» Men under tre dagar kunde de icke lösa gåtan.
Och om en kvinna i sin mans hus gör ett löfte, eller med ed förbinder sig till återhållsamhet i något stycke,
Asarja födde Heles, och Heles födde Eleasa.
Men Absalom sände ut hemliga budbärare till alla Israels stammar och lät säga: »När I hören basunen ljuda, så sägen: 'Nu har Absalom blivit konung i Hebron.'»
Herren kom såsom en fiende och fördärvade Israel, han fördärvade alla dess palats, han förstörde dess fästen; så hopade han över dottern Juda jämmer på jämmer.
Ingen som är född i äktenskapsbrott eller blodskam skall komma in i HERRENS församling; icke ens den som i tionde led är avkomling av en sådan skall komma in i HERRENS församling.
dit Gera jämte Naaman och Ahia förde bort dem: han födde Ussa och Ahihud.
Och HERREN sade till Samuel: »Huru länge tänker du sörja över Saul? Jag har ju förkastat honom, ty jag vill icke längre att han skall vara konung över Israel. Fyll ditt horn med olja och gå åstad jag vill sända dig till betlehemiten Isai, ty en av hans söner har jag utsett åt mig till konung.»
Och alla som bodde i Lydda och i Saron sågo honom; och de omvände sig till Herren.
De som då togo emot hans ort läto döpa sig; och så ökades församlingen på den dagen med vid pass tre tusen personer.
åt en gav han fem pund, åt en annan två och åt en tredje ett pund, åt var och en efter hans förmåga, och for utrikes.
När jag alltså vände mig till att jämföra vishet med oförnuft och dårskap -- ty vad kunna de människor göra, som komma efter konungen, annat än detsamma som man redan förut har gjort? --
Och deras barn talade till hälften asdoditiska -- ty judiska kunde de icke tala riktigt -- eller ock något av de andra folkens tungomål.
Ty tre äro de som vittna:
Han förde honom fram över landets höjder och lät honom äta av markens gröda; han lät honom suga honung ur hälleberget och olja ur den hårda klippan.
När de sedan gingo därifrån, bad men dem att de nästa sabbat skulle tala för dem om samma sak.
Och han åstundade att få fylla sin buk med de fröskidor som svinen åto; men ingen gav honom något.
Och HERREN gick förbi honom, där han stod, och utropade: »HERREN! HERREN! -- en Gud, barmhärtig och nådig, långmodig och stor i mildhet och trofasthet,
Och han sade till honom: »Stå upp och gå dina färde. Din tro har frälst dig.»
Därför har icke heller det förra förbundet blivit invigt utan blod.
Och jag, Johannes, var den som hörde och såg detta. Och när jag hade hört och sett det, föll jag ned för att tillbedja inför ängelns fötter, hans som visade mig detta.
Om däremot allenast få år återstå till jubelåret, så skall han räkna efter detta, sig till godo, och betala lösen för sig efter antalet av sina år.
Då sade han till mig: Gå; jag vill sända dig åstad långt bort till hedningarna.'»
Och de församlade sig till Jerusalem i tredje månaden av Asas femtonde regeringsår,
Ett mjukt svar stillar vrede, men ett hårt ord kommer harm åstad.
Ja, må din hand vara upplyft över dina ovänner, och må alla dina fiender bliva utrotade!
Och han sade till dem: »Jag har högeligen åstundat att äta detta påskalamm med eder, förrän mitt lidande begynner;
Ty lika visst som Jesus, såsom vi tro, har dött och har uppstått, lika visst skall ock Gud genom Jesus föra dem som äro avsomnade fram jämte honom.
Och när hon har funnit den, kallar hon tillhopa sina väninnor och grannkvinnor och säger: 'Glädjens med mig, ty jag har funnit den penning som jag hade tappat bort.'
honom som befaller solen, så går hon icke upp, och som sätter stjärnorna under försegling;
Och alla heliga gåvor som Israels barn giva såsom en gärd, vilken de bära fram till prästen, skola tillhöra denne;
Sedan kallade Abimelek Abraham till sig och sade till honom: »Vad har du gjort mot oss! Vari har jag försyndat mig mot dig, eftersom du har velat komma mig och mitt rike att begå en så stor synd? På otillbörligt sätt har du handlat mot mig.»
Ty jag vet att I efter min död skolen taga eder till, vad fördärvligt är, och vika av ifrån den väg som jag har bjudit eder gå; därför skall olycka träffa eder i kommande dagar, när I gören vad ont är i HERRENS ögon, så att I förtörnen honom genom edra händers verk.»
för honom som förvandlar klippan till en vattenrik sjö, hårda stenen till en vattenkälla.
Men dessa som stå efter mitt liv och vilja fördärva det, de skola fara ned i jordens djup.
Och Jesus begynte åter tala till dem i liknelser och sade:
att de skulle föra drottning Vasti, prydd med kunglig krona, inför konungen, för att han skulle låta folken och furstarna se hennes skönhet, ty hon var fager att skåda.
Ja, min boning skall vara hos dem, och jag skall vara deras Gud, och de skola vara mitt folk.
Ty se, de som hava vikit bort ifrån dig skola förgås; du förgör var och en som trolöst avfaller från dig.
Och du skall föra fram hans söner och sätta livklädnader på dem.
Och den överskrift som man hade satt upp över honom, för att angiva vad han var anklagad för, hade denna lydelse: »Judarnas konung.»
Han skulle ock bliva en fader för omskurna, nämligen för sådana som icke allenast äro omskurna, utan ock vandra i spåren av den tro som vår fader Abraham hade, medan han ännu var oomskuren.
