Vid tidsbeställningen får du veta hur snabbt du kommer att få vård.
Vanda centrum ligger i Dickursby.
Användarpanelen är öppen för alla som är intresserade av InfoFinland.
Du hittar mer information på HRT:s webbplats.
Rådgivning för ungafinska
Bostadsrättsbostad
Vilka hälsotjänster kan du använda?
På InfoFinlands sida Problematiska situationer i Helsingfors får du information om var i Helsingfors man kan få hjälp med barns och ungas problem, eller vid problem i familjen.
Om studeranden har ett annat modersmål än finska eller svenska och saknar tillräckliga språkkunskaper för gymnasiestudierna, kan hen söka till förberedande gymnasieutbildning (LUVA).
Senioruniversitetet (ikäihmisten yliopisto) är avsett för dem som har fyllt 60 år.
Det finska språket och den finländska kulturen och ekonomin utvecklades enormt under Finlands tid som en del av Ryssland.
Inga ytterligare begränsningar – Du får inte tillämpa lagliga begränsningar eller teknologiska metoder som juridiskt begränsar andra från att gör något som licensen tillåter.
På mötet kan man komma överens om hur situationen ska lösas.
Om du av någon anledning inte till exempel lyckas få en läkartid utanför arbetstiden, ska du komma överens med din chef om att du är borta och hur du ersätter din frånvaro.
En del av tjänsterna i Päihdelinkki finns även på svenska, engelska och ryska.
Kvällar och veckoslut är jourmottagningen centraliserad till större vårdenheter.
Rovala-institutets utbildning för invandrare
Lyft fram sådana färdigheter som behövs i uppgiften.
Läs mer på InfoFinlands sida Trafiken i Finland.
Om du har slutat använda preventivmedel, men en graviditet inte har börjat inom ett år, boka tid på hälsostationen eller hos en privat gynekolog.
En ung som inte är trygg i sitt eget hem kan kontakta Finlands Röda Kors De ungas skyddshus.
Som orsak för abort (abortti) räcker även att det med tanke på din livssituation skulle vara en alltför stor belastning att föda barnet eller att ta hand om det.
Vid mödrarådgivningen (äitiysneuvola) följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
Adjö.
Be om intyget av din arbetsgivare.
Om det är svårt eller omöjligt att bo i bostaden under reparationerna, har du rätt att säga upp hyresavtalet eller får nedsatt hyra.
Statsförvaltningens språkexaminafinska _ svenska
Även våld mot familjemedlemmarna är ett brott.
Du kan påvisa dina yrkeskunskaper med ett fristående yrkesprov.
Vanda och hela huvudstadsregionen har goda kollektivtrafikförbindelser.
registreringsintyget över uppehållsrätt för EU-medborgare (om du är EU-medborgare)
Assistenten kan hjälpa dig till exempel med att laga mat, handla, på din arbetsplats, i dina studier eller dina hobbyer.
Om du har din hemkommun i Esbo kan du utnyttja de offentliga hälsovårdstjänsterna.
En myndighet, till exempel en notaries publicus, måste verifiera överenskommelsen.
Webbplatsen betjänar även myndigheter i deras flerspråkiga informationsverksamhet.
företagsverksamheten är din huvudsyssla
Våld i hemmet
Anhållan om prövning av hinder mot äktenskapfinska _ svenska _ engelska
Då måste samhället ingripa i familjens situation.
Du kan även gå till en privat tandläkarmottagning.
Vårdbidrag för pensionstagare
Information om riksdagsvalfinska _ svenska _ engelska
Särskilt lönar det sig att utreda bostadens skick grundligt.
När du väntar barn
Dessutom används nationella läroplansgrunder och lokala läroplaner.
Om du har en bil måste du teckna en trafikförsäkring (liikennevakuutus).
Finland förlorade båda krigen, men Sovjetunionen ockuperade aldrig Finland.
Volontärarbetefinska
linkkiEures-portalen:
Dessa ordnas oftast i årskurs nio.
När du söker till ett universitet, får du i allmänhet poäng utifrån studentexamen och inträdesprovet.
hur många år du återbetalar lånet
linkkiFinska ortodoxa kyrkan:
Vilka tjänster ditt lands beskickning tillhandahåller beror på lagen i ditt hemland.
Arbetslagstiftningfinska _ svenska _ engelska
Meddela alltid
Också polisen kan undersöka orsaken till dödsfallet.
Integrationsrelaterade socialtjänster
På våren är det mycket svårt att bedöma isens bärkraft och då är det bäst att undvika att färdas på isen.
Tidsbeställning på vardagar.
Du kan även ringa kristelefonen om du är orolig för en närstående person.
I Esbo finns dessutom familjedagvårdare.
Registrering av uppehållsrätt för EU-medborgarefinska _ svenska _ engelska
Information om TE-byråns tjänster för invandrare finska _ svenska _ engelska
När föräldrarna skiljer sig ska de komma överens om underhållet av barnet samt om eventuellt underhållsbidrag (elatusapu).
Om ditt fostervatten går eller du har tätt återkommande smärtsamma värkar ska du ringa sjukhuset och fråga om det är dags att åka.
Om du inte har en bostad eller om du har bostäder på flera kommuners område är din hemkommun den kommun som du själv uppfattar som din hemkommun och som du har någon fast förbindelse till, till exempel genom familjeförhållanden eller arbetsplats.
Råd i frågor som rör familjen
Jämställdhet mellan män och kvinnor
I vissa fall kan du också få bostadstillägg, till exempel om du studerar på en avgiftsbelagd linje vid en folkhögskola och bor på läroanstaltens internat.
Be Fpa om mera information.
Det betyder att den som avlägger utbildningen får en arbetsplats hos arbetsgivaren.
Begravningsplatserfinska _ svenska _ engelska
Köp hållbara produkter.
Du måste betala avgiften samtidigt som du ansöker om fortsatt uppehållstillstånd.
Låt ögonläkaren undersöka dina ögon regelbundet så att eventuella ögonsjukdomar upptäcks i ett tidigt skede.
Efter att betänketiden gått ut ska du eller ni ansöka om slutlig äktenskapsskillnad inom ett halvt år.
Storleken på hyran varierar beroende på bostadens läge.
På vissa bibliotek ordnas även språkcaféer i det finska språket för invandrare.
tfn 0400 979 175
Friluftsområdenfinska _ svenska _ engelska
7–17-åringar har läroplikt (oppivelvollisuus), d.v.s. skyldighet att avlägga grundskolans (peruskoulu) lärokurs.
Du kan redogöra för hur du försörjer dig i Finland.
I Helsingfors finns många gymnasieskolor.
Finland är det viktigt att känna till de grundläggande reglerna som gäller i arbetslivet och det finländska samhället.
Du kan få hjälp med din rädsla till exempel vid polikliniken för förlossningsrädsla (synnytyspelkopoliklinikka).
Tänk på att arbete som freelancer eller företagare kan påverka din arbetslöshetsförsäkring.
Du kan också ansöka om många slags uppehållstillstånd och EU-registrering på internet i tjänsten Enter Finland.
I Esbo finns flera yrkes- och amatörteatrar.
Grundläggande utbildning
Barnet måste delta i förskoleundervisningen.
Information om företagshälsovårdenfinska _ svenska _ engelska
ditt utbildningsbehov
Offentliga hälsovårdstjänster tillhandahålls till exempel vid hälsostationer, tandkliniker, rådgivningsbyråer och sjukhus.
Arbets- och näringsbyrån väljer studerandena till den yrkesinriktade arbetskraftsutbildningen.
Magistraten fattar beslut om registrering av hemkommun.
I Helsingfors beslutas ärenden av stadsfullmäktige.
I början av året skickar staden en anmälan om läroplikt (oppivelvollisuusilmoitus) till hemmen.
I Finland fästs stor uppmärksamhet vid arbetssäkerhet.
Om du behöver akut tandläkarvård kvällstid eller under veckoslut, kan du kontakta Haartmanska sjukhuset i Helsingfors.
Du kan berätta vilka målsättningar du har med jobbsökningen eller vilken specialkompetens du besitter.
På webbplatsen för Suomen lakiopas får du information om vilka handlingar du behöver för bodelningen.
Om barnet inte är finsk medborgare måste han/hon ha uppehållstillstånd i Finland.
Tfn 075 7575 100
Gör videoklippet på något av de språk som används i Infobanken.
Mottagningscentralen betalar mottagningspenning till asylsökande.
Vi använder cookies
Jourmottagningen tar endast hand om barn med brådskande hjälpbehov.
I Helsingfors finns även ett muslimskt daghem vars verksamhetsspråk är arabiska.
Vilka möbler som ingår varierar.
Att ansöka om bostadsbidragfinska _ svenska _ engelska
Vetenskaplig fortbildning vid universitet
InfoFinland finansieras av staten och samarbetskommunerna.
Familjevård kan även ordnas i den vårdbehövandes eget hem.
Flyktingar kan be om hjälp och rådgivning i rättsliga frågor bland annat från flyktingrådgivningen r.f. eller från rättshjälpsbyråer.
Miessakit rf strävar efter att sörja för mäns välbefinnande och erbjuder sociala aktiviteter och stöd.
databehandling och datakommunikation
Närbiblioteken finns i Björkhagen, Kelviå, Lochteå samt Ullava kyrkby och Rahkonen.
Diskriminering på arbetsplatsen
Läs mer på InfoFinlands sida Brott.
Seniorernas tjänster, hemvårdfinska _ svenska
Om du är under 25 år, kontrollera tilläggsvillkoren för arbetsmarknadsstödet för unga på TE-tjänsternas webbplats.
Bokföring
Lagar och kollektivavtal reglerar exakt när tidsbundna anställningar får tillämpas.
Barnatillsyningsmännen ger även råd till föräldrar som ska skiljas.
I Finland gäller allemansrätten (jokamiehenoikeus).
Barns tandvård
Fråga om integration på svenska när din inledande kartläggning och integrationsplan görs.
Fråga vid socialbyrån om kommuntillägg betalas i din kommun.
Vi läser tillsammans i Vandafinska _ svenska _ engelska
Om du hemma vårdar en långtidssjuk, handikappad eller äldre familjemedlem kan din hemkommun betala stöd för närståendevård (omaishoidontuki) till dig.
Invandrarelever använder i huvudsak grundskolans och gymnasieskolans vanliga tjänster.
du kommer till Finland för att arbeta som tolk, lärare, sakkunnig eller idrottsdomare i högst tre månader utifrån en inbjudan eller ett avtal;
Du kan bo i bostadsrättsbostaden så länge du vill.
Undervisningsgruppen ska ha minst fyra elever.
Om du använder kollektivtrafiken ofta tjänar du på att ladda kortet med period.
linkkiFinlands Flyktinghjälp:
Som EU-medborgare kan du ansöka om studieplats vid en läroanstalt som är godkänd i Finland.
Det är viktigt att du har tillräckligt med kapital i startskedet.
Huvudstadsregionens gemensamma bibliotekstjänstfinska _ svenska _ engelska _ ryska _ somaliska _ persiska _ arabiska
Vaccinationer
I Vanda finns en delegation för mångkulturella frågor (monikulttuurisuusasiain neuvottelukunta) som lägger fram propositioner i ärenden som rör invandrare.
Engelsk-finskspråkigt daghemfinska _ engelska
Uppehållstillstånd på en ny grundfinska _ svenska _ engelska
Bolagsman i ett öppet bolag
Om din företagsverksamhet upphör, kan du ansöka om inkomstrelaterad dagpenning (ansiosidonnainen päiväraha) vid arbetslöshetskassan.
Du kan få arbetslöshetsstöd från och med det datum då du anmälde dig som arbetslös.
linkkiSkatteförvaltningen:
I särskilda fall kan barnet börja skolan senare.
Boka tid för vigseln hos magistraten eller tingsrätten i god tid före bröllopsdagen.
Du kan ansöka om moderskapspenning om du omfattas av den sociala tryggheten i Finland och varit sjukförsäkrad i Finland, ett annat EU- eller EES-land eller Schweiz oavbrutet i 180 dagar före det beräknade förslossningsdatumet.
Biträdet deltar i asylsamtalet efter sitt eget omdöme.
För registrering av en familjemedlem till en EU-medborgare krävs också att den person som är bosatt i Finland har tillräckliga medel för att försörja sig själv och sin familjemedlem som ska flytta till Finland.
För att du ska kunna få en hemkommun i Finland måste du flytta till och vara stadigvarande bosatt i Finland.
Evangelisk-lutherska församlingarfinska _ svenska _ engelska
linkkiStatens rättshjälpsbyrå:
Arbete och entreprenörskap
Målet är att stödja barnets utveckling och välbefinnande.
Hur sorteras avfall?
Om du tänker köpa en bostadsaktie, ta då även reda på vilka renoveringar bostadsaktiebolaget planerar och vad de kostar.
Om du vill ansöka om en hyresbostad, fyll i en ansökningsblankett för hyresbostad på Espoon Asunnot Oy:s webbplats.
ni har gemensamma barn eller
Utkomststöd kan du få om du inte lyckas få tillräckliga inkomster genom eget arbete, andras omsorg eller på något annat sätt.
Du kan ansöka om en delägarbostad med en ansökan riktad till bostadens byggherre.
Serviceboende är en boendeform avsedd för sådana personer som behöver kontinuerlig hjälp men inte är i behov av anstaltsvård.
Du kan låta utföra ändringsarbeten i ditt hem som underlättar boendet.
Ungdomsgårdarfinska _ svenska _ engelska
Med sökmotorn kan du kontrollera var och när du kan avlägga examen.
linkkiUtbildningsstyrelsen:
Arbetstagaren kan få ersättning vid ett olycksfall.
Mer information får du till exempel på Väestöliittos webbplats eller webbplatsen för kyrkans familjerådgivningscentral.
Öppna yrkeshögskolor
På stadens webbplats finns även en länk till Evenemangskalendern med daglig information om stadens kultur- och motionsevenemang.
Du kan även beställa skattekortet via Skatteförvaltningens telefontjänst:
Ditt födelseår avgör i vilken ålder du kan få arbetspension.
Arbetstiden ska följa arbetslagstiftningen och kollektivavtalet.
Adress: Sörnäsgatan 1
Penningunderstöd för utländska forskarefinska _ svenska _ engelska
Läs mer: Högskoleutbildning
När du vill flytta behöver du inte sälja bostaden.
Du kan också lämna initiativ och ställa frågor samt kommentera ärenden på finska och på svenska.
Motion.
Hyresvärden ska meddela hyresgästen om hävandet.
P-EU-tillstånd gäller tills vidare.
legitimation (till exempel pass)
I Finland råder också yttrandefrihet.
Om man redan behärskar de färdigheter som krävs för examen, kan man också avlägga yrkesexamen eller specialyrkesexamen som yrkesprov.
Minimiarbetstiden är vanligtvis 18 timmar i veckan.
Samtalen är konfidentiella.
Rätten till en hemkommun i Finland bestäms enligt hemkommunslagen.
Val av förlossningssjukhusfinska _ svenska _ engelska
tfn 016 322 8091 eller tfn 016 322 8014
Hur ansöker man om en bostadsrättsbostad?
Om du flyttar ditt stadigvarande boende till Esbo, ska du registrera dig som invånare i kommunen.
Polisen utfärdar identitetskort.
Läs mer: Bibliotek
Avsikten är att fadern tar hand om barnet.
Föräldrarna kan hjälpa ledarna att utarbeta planen.
Om din arbetsgivare är finländare eller om din utländska arbetsgivare har en arbetsplats i Finland, betalar du skatt i Finland.
Hyresgästen har rätt att göra detta, om bostadens egentliga hyresvärd godkänner detta.
Mer information om motionsrutterna, rastplatser, möjligheter till fiske och båtliv samt exempelvis fågeltorn i Karleby finns på stadens webbplats.
tfn (09) 839 22133
Tjänsten är kostnadsfri.
Om du är medborgare i något av de nordiska länderna, ett EU-land, ett EES-land eller i Schweiz och kommer till Finland för att arbeta, behöver du inget uppehållstillstånd.
Läs mer: Fritid i Esbo
I den finländska kulturen följs dock fortfarande många kristna seder.
1918 Inbördeskrig mellan röda och vita
Du kan skriva ut blanketten på Migrationsverkets webbplats.
Om ett barn blir akut sjukt, ska du ta kontakt med hälsostationen eller jourmottagningen.
Statsförvaltningens språkexamen om kunskaper i finska och svenska
Allmänt bostadsbidragfinska _ svenska _ engelska
De flesta webbkurser är på finska eller svenska, men det finns även andra alternativ:
Om arbetsgivaren säger upp en arbetstagare måste arbetsgivaren ange orsaken till detta.
I Finland finns många föreningar för invandrare.
Helsingfors är Finlands administrativa centrum: där sammanträder Finlands riksdag och där finns ministerierna.
Även om Helsingfors växte snabbt, var Esbo ännu länge en fridfull landssocken.
Besök läkaren
När du registrerar ditt företag för första gången ska du fylla i en etableringsanmälan och skicka in erforderliga bilagor.
I Esbo finns många olika hotell där man kan bo tillfälligt.
Kompetenscentret Stadin osaamiskeskus (Stadin osaamiskeskus) förbereder invandrare för arbetsmarknaden och hjälper dem att hitta ett jobb eller en praktikplats.
Du kan söka en jurist till exempel på Finlands advokatförbunds webbplats, via tjänsten Etsi asianajaja.
Använd inte vatten.
Det är också viktigt att du bekantar dig med finländare och arbetslivet i Finland redan under studietiden.
avsluta inte samtalet förrän du får lov.
Även om du väljer integrationsutbildning på svenska lönar det sig för dig att i något skede även lära dig finska.
Begravningsbyråer hjälper med de praktiska arrangemangen vid en begravning.
Kompetenscentret för integration av invandrare stöder arbete som främjar integrationen av invandrare lokalt, regionalt och riksomfattande.
Vid tidsbeställningen bedöms vilken slags vård barnet behöver.
Du kan till exempel ta vilket som helst namn som du har haft tidigare.
du har rätt att använda arbets- och näringsbyråns tjänster.
Du kan även besöka FPA:s kontor.
Mer information hittar du på InfoFinlands sida Finska och svenska språket.
Friluftsområdenfinska
Brådskande ärenden är till exempel bihåleinflammation, ögoninfektion, ryggvärk, en lindrig urinvägsinfektion, en vaginal infektion eller eksem.
annan orsak
Vanligtvis börjar förskoleundervisningen det år då barnet fyller sex år.
Barnets officiella adress påverkar också till exempel FPA:s bostadsbidrag.
Sambo med en finsk medborgare
svåra livssituationer
Du kan få:
Om du vill läsa finska eller svenska, läs mer på InfoFinlands sida Finska och svenska språket.
specialyrkesexamina.
Om den egna hälsostationen eller det egna sjukhuset inte kan ge patienten vård inom utsatt tid måste de ordna möjlighet för patienten att få vård på ett annat ställe.
Flyttanmälan ska alltid göras till magistraten (maistraatti).
Om du kommer från ett annat EU-land kan du i vissa fall utnyttja de försäkringsperioder som du har ackumulerat i andra EU-länder.
Om du får mer lön än vad du uppgett, överskrids din inkomstgräns.
Arbetsmarknadsstödfinska _ svenska _ engelska
Under Stora nordiska kriget år 1710 föll två tredjedelar av Helsingfors befolkning offer till pesten.
FöretagsFinland (via webbplatsen och per telefon)
Broschyren Jobba i Finland(pdf, 5,51 MB)finska _ svenska _ engelska _ ryska _ estniska _ franska _ polska
Biskopsbron 9 B
Sambo till en person som fått internationellt skyddfinska _ svenska _ engelska
Ett barn eller barnbarn under 21 år som är beroende av din sambo för sin försörjning
Vem kan ställa upp som kandidat?
Detta innebär att du på förhand betalar ett penningbelopp som motsvarar några månaders hyra till hyresvärden.
Familjerådgivningen betjänar invånarna i Grankulla.
Om du vill ansöka om finskt medborgarskap (kansalaisuus) kan du påvisa att du har tillräckliga kunskaper i finska eller svenska genom att avlägga den muntliga och skriftliga delen av en allmän språkexamen minst på nivå 3.
humanistiska och konstnärliga områden
De strävar efter att förbättra dessa minoriteters ställning i samhället.
Han eller hon kan således inte hjälpa dig med annat.
Seniorrådgivningenfinska _ svenska _ engelska
Den ordnas i daghemmens förskolegrupper.
Tjänsten kan också användas av andra invandrare som behöver tillfällig rådgivning i specialfrågor som rör integration.
Information om vård av drogproblemfinska _ svenska _ engelska
Dessutom ska ditt barn ha en finländsk personbeteckning.
Statsborgen kan utgöra högst 20 procent av lånet och högst 50 000 euro.
Fråga din arbetsgivare som det ordnas undervisning i det finska språket på din arbetsplats.
Boendeguide för ungafinska
Vid arbetarinstitutet kan vem som helst studera.
Återvinningsstationerfinska _ svenska _ engelska
Utöver skatt betalar arbetsgivaren försäkringspremier på din lön i händelse av arbetslöshet eller sjukdom.
Alla länder har inte en beskickning i Finland.
modern har en finsk personbeteckning.
Mer information om att köpa en egen bostad får du på banken eller hos fastighetsförmedlare.
Muslimernas gravkvarterfinska
Som studerande betalar du själv vårdkostnaderna om du insjuknar i Finland.
Också Helsingfors församlingar har klubbverksamhet.
nyårsdagen 1.1
Vid Karleby finska gymnasium anordnas undervisning i finska som andraspråk för invandrare invandrare.
mån kl. 9–16 utan tidsbeställning
Diskriminering är ett brott.
Sommaruniversitets kurser är avgiftsbelagda för deltagarna.
Information om gymnasiestudierfinska _ svenska _ engelska
Lämna eller posta blanketten till den dagvårdsenhet där du i första hand söker plats.
Äktenskap mellan följande nära släktingar är förbjudet:
Observera att utländska handlingar ska vara legaliserade.
Vuxenutbildningsinstitutet ordnar även kurser för invandrare.
Gör flyttanmälan senast inom en vecka från din flyttningsdag.
Karleby stads blankett för ansökan om hyresbostad kan fyllas i och skickas in på nätet.
Yrkesutbildning efter gymnasiet
studerande
Vissa spermiedödande medel kan köpas receptfritt på apotek.
Om du till exempel har bokat tid hos en myndighet eller läkaren är det speciellt viktigt att du är på plats i tid.
Vanligen består ett hushåll av ett äkta par, sambor eller en familj.
Studier i finska språket på Internetfinska _ engelska
Hindersprövningen görs på magistraten (maistraatti).
Även om du har kommit lagligt till Finland kan din vistelse i landet bli illegal till exempel om du stannar kvar i landet fastän du inte beviljas ett uppehållstillstånd eller om ditt visum eller uppehållstillstånd har gått ut.
Till exempel ska lokaler där man säljer livsmedel eller idkar skönhetsvård kontrolleras och tillstånd sökas hos kommunens hälsomyndighet innan lokalerna tas i bruk.
Om du till exempel har en krävande hobby eller är sjuk en lång tid kan du avlägga gymnasiet som distansstudier.
Barnet kan få minst 20 timmar småbarnspedagogik i veckan eller mer om föräldrarna arbetar eller struderar.
bostadens storlek
Jourmottagningarfinska _ svenska _ engelska
Ansökan till yrkesutbildning
Skattenummer
linkkiFlyktingrådgivningen r.f.:
linkkiMellersta Österbottens folkhögskola:
Ingen får behandlas annorlunda till exempel på grund av kön, ålder, religion eller handikapp.
Det finns olika CV-mallar.
Här kan du hämta ett skattekort och ett inom byggbranschen obligatoriskt skattenummer.
Förlossningen
Du kan söka information om rutterna i reseplanerartjänsten (Reittiopas).
Den första finskspråkiga ABC-boken (Aapinen) ges ut i Finland
Under den förberedande undervisningen studerar barnet eller den unga finska och några läroämnen.
Att köra bil under alkoholpåverkan är förbjudet enligt lag och det kan ge ett hårt straff.
Ersättningen kan vara en ersättning av sjukvårdskostnader och inkomstbortfall i form av dagpenning, olycksfallspension, ersättning för den skada som olyckan har orsakat, rehabilitering eller vid dödsfall familjepension till de anhöriga.
I Karlebynejden erbjuds olika inkvarteringsalternativ.
Åldringar kan använda tjänsterna vid de vanliga hälsostationerna.
I Finland har barn rätt till särskilt skydd och särskild omsorg.
Vid problem med din mentala hälsa ska du i första hand kontakta din egen hälsostation eller företagshälsovårdens mottagning.
Om ditt land har tillträtt Haagkonventionen ska du begära om ett så kallat Apostille-intyg för din handling.
Jag hittar inte en förmånlig hyresbostad.
Uppfostring av barn i Finland(pdf, 8,08 Mt)finska _ engelska _ ryska _ somaliska _ kurdiska _ albanska _ burmesiska
Helsingfors evenemangskalenderfinska
När du vill starta ett företag ska du fundera noga på om du har en bra affärsidé.
Om du har kommit till Finland som kvotflykting, kan Migrationsverket ersätta kostnaderna för en familjemedlems inresa.
NEJ: glasföremål, glaskärl, speglar, porslin
Telefontjänst: 0295 020 500
Anmäla födelsen av ditt barn till myndigheterna i ditt hemland om barnet föds i Finland
Läs mer om arbetslöshetskassan på InfoFinlands sida Fackförbund.
linkkiYrkesutövarnas och företagarnas arbetslöshetskassa:
Om samborna förvärvar egendom tillsammans ska båda parterna antecknas som köpare och alla kvitton sparas.
Läroavtalsplatsen kan också vara din nuvarande arbetsplats.
Om du inte har en sådan handling, kan dina fingeravtryck jämföras med de fingeravtryck som lagrats i uppehållstillståndskortet eller uppehållskortet.
Karleby hamn ligger i stadsdelen Yxpila och är en av Finlands mest trafikerade godshamnar.
Kom ihåg att företagande även medför risker.
Genom att betala en bostadsrättsavgift, som är 15 procent av bostadens anskaffningspris, och därefter varje månad ett rimligt bruksvederlag får man rätt att förvalta över bostaden precis som om den vore en ägarbostad.
Företagarkurser
Telefonrådgivning: 0295 666 842
Arvsskatt
Flyktingar kan även kontakta Esbo stads invandrartjänster (Maahanmuuttajapalvelut).
Företagare i Esbo får även hjälp av Företagarna i Esbo rf.
I Finland finns 40 nationalparker.
När flyktingarna anländer till Finland kommer en anställd från röda korset till flygplatsen och tar emot dem.
Vissa museers samlingar kan du även bekanta dig med på internet.
Diskrimineringsombudsmannen kan ge anvisningar, råd och rekommendationer samt hjälpa parterna att åstadkomma förlikning i diskrimineringsfall.
Vailla vakinaista asuntoa ry har ett nattcafé, Kalkkers, som erbjuder bostadslösa en varm plats på natten från höst till vår.
Biblioteket producerar även läroböcker för synskadade skolelevers och studerandes behov.
Kondomer säljs också till exempel i mataffärer.
Migrationsverket beslutar om du får uppehållstillstånd eller inte.
Om du och din granne har en konflikt som ni inte klarar av att själva lösa, kan ni be om hjälp vid grannmedlingscentret Naapuruussovittelun keskus eller hos disponenten.
Graviditet kan också förhindras med spermiedödande medel, till exempel p-skum (emätinvaahto) eller slidpiller (emätinpuikko), men de är inte särskilt effektiva.
Läs mer: Studier som hobby
Webbkurs med många hjälpspråksvenska _ engelska _ ryska _ franska _ spanska _ kinesiska _ tyska _ portugisiska
Familjeplanering
Anvisningar om eftermiddagsverksamhetens klientavgiftfinska _ ryska _ somaliska _ arabiska
På museiförbundets sidor hittar du mer information om dagar med fritt inträde.
Sådana hjälpmedel är till exempel datorer och tilläggsutrustning till datorer.
Kontrollera ersättningen i ditt kollektivavtal.
linkkiRegionförvaltningsverket:
Ansök om fortsatt uppehållstillstånd elektroniskt i tjänsten Enter Finland eller på Migrationsverkets tjänsteställe.
Både myndigheter och vanliga människor deltar i flaggdagarna.
Magistraten registrerar dina uppgifter i det finska befolkningsdatasystemet.
Barnet behåller sitt tidigare efternamn när föräldrarna skiljer sig.
börjar det år då barnet fyller 7 år
VALMA-utbildningen räcker ungefär ett läsår.
I arbetslivet syns religionens inflytande i de många lediga dagarna som anställda får.
linkkiKarleby kyrkliga samfällighet:
Du behöver inte tillstånd av dina föräldrar för receptet.
Du betalar avgiften när du lämnar in din tillståndsansökan.
Flygplatsen finns i Kronoby på endast 22 kilometers avstånd från Karleby centrum.
Information om tandvårdenfinska _ svenska _ engelska
Sök tandläkarefinska
Grankulla hälsostation
Motiverade skäl för förlängning av visum kan till exempel vara:
Kurserna är avgiftsbelagda och de ordnas både dag- och kvällstid.
Tolkning för en handikappad är inte det samma som språktolkning.
Förmånliga utlandssamtalfinska _ svenska _ engelska
Självständiga språkanvändare
Ämnen som behandlas på kurserna är till exempel utarbetande av en affärsverksamhetsplan, startande av företagsverksamhet, bokföring, företagsbeskattning, juridiska frågor, marknadsföring, försäljning och kundtjänst.
Avgiften är ca 15 procent av bostadens pris.
Delta i tävlingen med ditt eget videoklipp!
Då är du återflyttare (paluumuuttaja).
Information om TE-byråns tjänster hittar du på InfoFinlands sida Om du blir arbetslös.
Närmare kontaktuppgifter finns på Esbo stads webbplats.
Om du på grund av skada eller sjukdom inte kan arbeta kan du få invalidpension (työkyvyttömyyseläke).
Den finansieras med skattemedel och är därför förmånligare för familjerna.
När äktenskapets lagliga villkor uppfylls kan ett par gifta sig.
När du går till magistraten ska du ta med dig
I Finland äter man lunch tidigare än i många andra länder.
linkkiTjänstemannacentralorganisationen STTK:
linkkiFinland-Samfundet:
Därefter övergår eleven till en vanlig klass.
På många metrostationer kan du parkera din bil gratis för att fortsätta resan med kollektivtrafiken.
Finland som en del av Sverige och Ryssland
Mer information om anmälan får du på Utbildningsstyrelsens (Opetushallitus) webbplats.
Att ansöka om partiell sjukdagpenningfinska _ svenska _ engelska
Körkort
Utlänningar som bor stadigvarande i Finland och som har fyllt 18 år har rätt att rösta i kommunalval.
Tidsbokning och rådgivningfinska _ svenska _ engelska
Karlebystödfinska _ svenska
Ofta ingår rättsskyddsförsäkringen i hemförsäkringen.
På motionsslingorna kan man springa på somrarna och åka skidor på vintrarna.
Du kan söka till dessa utbildningar i den kontinuerliga ansökan året om eller i den gemensamma ansökan till andra stadiet.
Vid behov kan du försöka förhandla om att avsluta hyresavtalet tidigare.
Betalningen av utkomststöd påverkas av alla dina inkomster och tillgångar.
Mödrahemmets tjänster är avsedda för personer som har hemkommun i Finland.
nattetid kl. 22–8
Badhuset/simhallen Vesihiisi
Munhälsovårdenfinska _ svenska
Läs mer om Inkomstregistret och om att anmäla löner på Inkomstregistrets webbplats.
Vid hälsopunkten Daalia ges vägledning och rådgivning för personer över 65 år om diet, motion och livsstil.
Studiebostäderfinska _ engelska
Information om Finlands historiaengelska _ ryska _ franska _ spanska _ tyska _ portugisiska
identitetsbevis (till exempel pass)
Du får studiehandboken till exempel på bibliotek eller Vandainfo samt i elektroniskt format på Vanda stads webbplats.
Det grundläggande utkomststödet täcker även utgifter för hobby- och rekreationsverksamhet, avgifterna för barndagvård och för skolbarns morgon- och eftermiddagsverksamhet samt nödvändiga kostnader för flytt.
Arbetsgivaren har skyldighet att:
Du ska söka med en separat ansökan t.ex.
Uppsägningstid
En del privata läkarstationer erbjuder denna tjänst. Ett hembesök av en privatläkare är dock dyrt.
Jämför olika mäklarbyråers priser på förhand.
Mer information om den förberedande undervisningen för invandrare får du av stadens undervisningstjänster.
Yles radiokanal Mondo erbjuder radioprogram på engelska och många andra språk.
Uppehållstillstånd för studerande beviljas högst för två år i taget.
Gränskontrollmyndigheten eller polisen registrerar dig som asylsökande, antecknar uppgifter om dig och tar dina fingeravtryck.
Flerfaldigt medborgarskap
Man kan resa nästan över allt i Finland med tåg eller buss.
Barns och ungas problem
studieplats
Är jag offer för människohandel?
Föreningen för bostadslösafinska _ engelska
Faderskapet kan erkänns redan under graviditeten vid mödrarådgivningsbyrån eller efter barnets födelse hos barnatillsyningsmannen i den egna kommunen.
Läs mer: Hälsovårdstjänster i Finland.
Flyktingar och asylsökande samt andra utlänningar kan söka hjälp och råd i frågor kring uppehållstillståndet hos Flyktingrådgivningen rf.
När du söker asyl utreder Migrationsverket samtidigt om du kan få uppehållstillstånd på någon annan grund.
Idrottstjänsterfinska _ svenska _ engelska
Kontrollera regelbundet att vattenledningarna i ditt hem inte läcker och att det inte rinner ut vatten från hushållsapparaterna på golvet.
Du kan hämta en personbeteckning och samtidigt registrera ditt tillfälliga boende i den närmaste magistraten (maistraatti) eller skattebyrån (verotoimisto).
Då du kommer till sjukhuset ska du använda centralsjukhusets huvudingång kl. 7–20 och övriga tider bör du använda den gemensamma jourens/poliklinikens dörr.
Mer information får du via tjänsten Helsingforsregionen.fi.
Förskoleundervisningen börjar i augusti och ansökningstiden är i januari.
Bostäder för bostadslösafinska
Information om skyddshem och mödrahemfinska
Om du inte får hjälp av din förman ska du ta kontakt med arbetsplatsens arbetarskyddsfullmäktige (työsuojeluvaltuutettuu) eller förtroendeman (luottamusmies).
Det är inte tillrådligt att säga upp hemförsäkringen under tiden då du bor i bostaden.
När man talar om lön avser man oftast bruttolönen (bruttopalkka) från vilken skatter och personalbikostnader dras av.
De annonseras inte ut öppet, utan arbetsgivarna söker arbetstagare via sina egna nätverk.
Parförhållandet registreras på magistraten.
Du hittar information om arbetstagarens rättigheter och skyldigheter i Finland på InfoFinlands sida Arbetstagarens rättigheter och skyldigheter.
Dessutom erbjuder även privata musikskolor och -institut undervisning.
Vissa inträdesprov omfattar förhandsuppgifter.
Skattefinska _ svenska _ engelska
Om du har hemkommun i Finland.har du rätt att få dessa undersökningar gjorda.
Du kan ansöka om stöd för närståendevård hos socialbyrån i din hemkommun.
Om du misstänker att barnets hälsa eller säkerhet äventyras när barnet träffar den andra föräldern ska du meddela detta till socialmyndigheter.
finska 029 497 000
Observera att tull- och skattefriheten för flyttsaker inte gäller alkohol eller tobaksprodukter.
Mer information om jämställdhet hittar du på InfoFinlands sida Jämställdhet och likabehandling.
Tandvårdens jourmottagning kvällar och veckoslutfinska _ svenska _ engelska
Är du studerande lönar det sig att ansöka om en studentbostad då dessa vanligen är förmånligare än andra hyresbostäder.
Mannerheims barnskyddsförbund MLL
Om du planerar adoption inom familjen ska du kontakta socialbyrån i din hemkommun.
om förlossningen kan utgöra en risk för din hälsa
Rådgivning för att motarbeta diskriminering
Området hade en direkt förbindelse till Helsingfors.
Stadslotsen har jour i områdets bibliotek vissa veckodagar och klockslag.
Fyll ansökan i tjänsten Studieinfo.fi.
Bostäder säljs av privatpersoner, fastighetsförmedlingar och byggherrar.
På Väestöliittos webbplats hittar du information om olika preventivmedel.
Läroanstalten kan kontrollera att du har tillräckliga språkkunskaper för studierna.
Basfakta
Det betjänar invandrare som är bosatta i Rovaniemi och annorstädes i Lappland.
Du hittar urvalet av språk i tjänsten i menyn uppe på sidan.
Du kan lämna in ansökan om skilsmässa till tingsrätten i din egen eller din makas/makes hemkommun.
Läs mer:
Rehabiliteringspenningfinska _ svenska _ engelska
möbler och andra husgeråd
Hur ansöker jag?
Lån som beviljas av banker eller Finnvera är vanliga finansieringskällor för många nya företagare.
Du ska besöka tjänstestället inom tre månader efter att ha gjort ansökan.
– Om du vill kan du även lista dina publikationer eller arbetsprov.
Dessutom ska du ha hemkommun i Finland den 51:a dagen före valdagen.
Om du inte är medborgare i något av Europeiska unionens medlemsländer, ett EES-land eller i Schweiz och vill driva ett företag i Finland, behöver du ett uppehållstillstånd för företagare.
Om du ska utföra säsongsarbete i Finland behöver du ett säsongsarbetstillstånd.
Mellersta Österbottens och Österbottens rättshjälpsbyrå
Läs mer: Barn vid skilsmässa
Du får mer information om att legalisera officiella handlingar vid magistraten eller beskickningen för ditt eget land i Finland.
Senare kan du köpa hela bostaden så att den blir helt och hållet din egen.
Vem kan få en bostadsrättsbostad?
Information för utvecklingsstörda och anhörigafinska
Största delen av verksamheten på ungdomsgårdarna är gratis.
Det är avgiftsfritt.
Om du har en hemförsäkring, och din bostad blir skadad till exempel vid en brand eller till följd av en vattenskada, kontakta då genast ditt försäkringsbolag.
Vi har samlat kontaktuppgifter till myndigheterna på InfoFinlands sida Ring och fråga om råd.
Om du ämnar flytta utomlands från Finland för två år, till exempel på grund av arbete eller studier, kan du ansöka hos Migrationsverket om att ditt uppehållstillstånd inte återkallas.
Detta måste du emellertid alltid komma överens om med hyresvärden.
linkkiMellersta Österbottens sommaruniversitet:
Religionsfrihet och religionsutövande i Finland
Efter grundskolan (peruskoulu), d.v.s. efter grundstadiet fortsätter studerandena till läroanstalter på andra stadiet (toisen asteen oppilaitos).
Tfn (09) 8789 1344
