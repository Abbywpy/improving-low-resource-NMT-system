Gör ansökan inom tre månader efter datumet för inresa.
En del tolkcentraler har jour på veckoslut samt kvällar och nätter.
kan den ena sambon inte få änkepension om den andra sambon dör.
Fundera också på om du har tillräckliga yrkeskunskaper och erfarenhet.
Karleby verksamhetsställe
transporttjänster
Använd inte elapparater som är i dåligt skick eller vars sladd är trasig.
Nuortenkatu 11
Läs mer på InfoFinlands sida Tjänster för handikappade.
Om du kommer som flykting till Finland ska du komma överens om en hälsokontroll med Utlänningsbyrån.
Ansvarsområdena för arbetarskydd ger både arbetstagare och arbetsgivare råd i frågor som gäller arbetets säkerhet och hälsa samt i frågor som rör anställningsvillkor.
är fadern förpliktad att delta i underhåll av barnet
Kvotflyktingar
Faderskapsledighet
Handläggning av ansökan om registrering av uppehållsrätt är avgiftsbelagd.
har det uppehållstillstånd (oleskelulupa) som krävs och
_ holländska _ kroatiska _ rumänska _ ungerska _ japanska _ italienska
Myndigheter som utfärdar Apostilleintyg finns i alla länder som är anslutna till Haagkonventionen.
Barnen har ofta en och samma lärare under de sex första skolåren.
FPA:s kunder är alla personer som bor i Finland och utomlands och som omfattas av socialskyddet i Finland.
Om det till exempel anges i hyresavtalet att det är förbjudet att röka i bostaden, kan du inte röka i ditt hem.
Om äktenskapet till exempel har varat under fem år delas egendomen inte nödvändigtvis jämnt.
Barnbidraget för det första barnet uppgår till cirka 100 euro per månad.
Jorvs sjukhus
I Finland visas filmerna oftast på originalspråket.
Arbets- och näringsbyråerna och kommunerna tillhandahåller invandrarrådgivning.
Behovsprövad rehabiliteringfinska _ svenska
Om du inte tar emot platsen i tid, förlorar du den.
När du inleder företagsverksamheten har du många skyldigheter, bland annat ska du registrera företaget och ordna beskattning och bokföring.
Om du redan är i Finland och får ett negativt beslut om uppehållstillstånd från Migrationsverket (Maahanmuuttovirasto), måste du antingen lämna Finland eller överklaga beslutet.
Till ansökan om uppehållstillstånd för arbetstagare ska du bifoga blanketten TEM054 som din arbetsgivare fyller i och undertecknar.
Till exempel på Helsingfors stads webbplats finns en färdig blankett, ett responssystem (palautejärjestelmä).
Om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
När ni kräver bodelning förordnar tingsrätten en bodelningsman som delar egendomen.
Sanduddsgatan 5 B
Du hittar kontaktuppgifterna på Sopu-arbetets webbplats.
Arbetstagare, företagare, studerande, flykting, asylsökande eller en familjemedlem till en person bosatt i Finland hittar information speciellt om sin egen situation på dessa sidor i Infobanken.
Du får hjälp med spelproblem vid A-kliniker (A-klinikka), mentalvårdsbyråer (mielenterveystoimisto) och hälsovårdscentralen (terveyskeskus).
Om du blir bostadslös, kontakta Esbo stads verksamhetsställe för vuxensocialarbete.
Tjänsterna och priserna i olika flyttfirmor kan variera stort och därför lönar det sig att jämföra.
I Vanda finns 10 bibliotek (kirjasto) och två bokbussar (kirjastoauto).
Infomötena är avgiftsfria.
Det kan vara fördelaktigt att kunna svenska när du söker jobb.
Startpenning
ensamboende eller
Stöd för skolresor
I Finland kan du avbryta en graviditet i tidigt skede i följande fall:
Om dina studier fortsätter men uppehållstillståndet håller på att gå ut ska du ansöka om fortsatt uppehållstillstånd.
Information om priser på sålda bostäderfinska _ svenska
Mun- och tandhälsovårdenfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster:
När din examensnivå har jämställts med en finländsk högskoleexamen, kan du söka till uppgifter som kräver den nivå på högskoleexamen som du har.
Skriv alltid ett skriftligt anställningsavtal innan du börjar på ett nytt jobb.
I de allra nordligaste delarna av Finland går solen inte alls ner i början av sommaren.
någon hotar dig eller din familj med våld
Information om boendefinska _ engelska
Barnen äter en varm måltid i skolan.
Mer information om juristtjänster och rättshjälp hittar du på InfoFinlands sida Behöver du en jurist?.
Heminkvarteringengelska _ franska _ spanska _ kinesiska _ tyska _ portugisiska _ italienska
När du ansöker om startpeng undersöker TE-byrån om företagandet är ett lämpligt alternativ för dig.
Finländare väntar vanligtvis att samtalspartnern har sagt sitt innan de själva tar till ordet.
linkkiFörbundet för Steinerpedagogik:
Om du inte förstår finska eller det finska teckenspråket kan du också behöva en annan tolk.
Du kan söka olika föreningar i patent- och registerstyrelsens tjänst Föreningsregistret.
I arbetsavtalet fastställs arbetsuppgifterna och lönen samt andra förmåner och villkor.
Om din arbetserfarenhet i Finland är kort eller om din finska ännu inte är så bra, kan frivilligarbete vara ett bra sätt att få fotfäste i arbetslivet och förbättra språkkunskaperna.
Boende i bostadsrättsbostad
(Det är bra att veta att stadigvarande boende definieras på olika sätt i olika lagar.
Under prövotiden kan arbetstagaren och arbetsgivaren häva arbetsavtalet utan uppsägningstid.
Tfn 045 134 1711
Prästgårdsgränden 5
Läroplikten upphör när barnet har fullgjort hela lärokursen för den grundläggande utbildningen eller det har förflutit tio år sedan läroplikten började.
Företagare måste inte ordna företagshälsovård för sig själv, men däremot måste de ordna det för sina anställda.
Om du vill att en mäklare söker en lämplig hyresbostad åt dig, ska du ingå ett skriftligt uppdragsavtal (toimeksiantosopimus) med mäklaren.
Guide om att grunda ett företagfinska _ engelska _ kinesiska
linkkiEvangelisk-lutherska kyrkan i Finland:
Bostadslån
Om du upprepade gånger bryter mot husets ordningsregler har hyresvärden rätt att häva hyresavtalet.
Den som är en enskild näringsidkare beskattas på så sätt att alla inkomster som återstår efter att man har dragit av kostnaderna för företagsverksamheten är beskattningsbara inkomster.
Tillstånet kan dras tillbaka om du permanent flyttar från Finland, uppehåller dig utomlands kontinuerligt i minst två år eller har lämnar felaktiga uppgifter då du ansökt om tillståndet.
Detta är det bra att beakta när du väljer företagsform.
Gravplats
De flesta jobben är dolda jobb.
För vilka studier kan man få arbetslöshetsförmån?
Kontrollera detta med din arbetsgivare.
Nattcentret Kalkkersfinska
Både offret och förövaren kan få hjälp.
Finska medborgare kan i Finland dömas för brott som begåtts utomlands.
Till exempel utbytesstuderande får inte finskt studiestöd.
Du ska också ha en giltig trafikförsäkring (liikennevakuutus) för din bil i Finland.
Vardera maken ansvarar ensam för den skuld som de har tagit före äktenskapet eller under det.
Finlands historia är en berättelse om handelsvägar, möten mellan kulturer och livet intill stora grannar.
Undervisning i den egna religionenfinska
Brådskande psykiatrisk sjukvård ges på jourenheter vid psykiatriska sjukhus.
FöretagsFinland
Tfn (09) 622 4322
Stöd och handledning för ungafinska _ engelska
Flerspråkiga biblioteket
Närskolan är oftast den skola som ligger närmast barnets hem.
Du kan också köpa avgiftsbelagda kanaler.
Du måste ha med ett ID-kort när du röstar.
Fråga mer på din hälsostation.
Om du vistas i Finland i mer än sex månader, ska du i allmänhet betala skatt på din lön till Finland.
När du ansöker om startpenning utreder arbets- och näringsbyrån om företagande är ett lämpligt alternativ för dig.
För att kunna ansöka om en hyresbostad hos staden, måste du ha uppehållstillstånd för minst ett år.
Information om kurser i skidåkning, om att hyra skidor och om skidspår finns till exempel på Suomen Latu ry:s webbplats på finska.
Förberedande utbildning inför yrkesutbildning
Finest sänder radioprogram på estniska.
Experterna där hjälper dig att utveckla affärsidén. Du får hjälp med att utarbeta preliminära marknadsundersökningar, lönsamhetskalkyler och en kartläggning om tillgången till finansiering.
Olika instanser anordnar företagarkurser och informationsmöten som man har mycket nytta av om man vill starta ett företag.
Begäran om prövning kan ställas på vilken magistrat som helst.
Tfn 016 3222 570.
Du ska ta pillret så snart som möjligt efter samlaget, i regel senast inom 72 timmar.
Karlebygatan 74
Dagvårdsavgifterfinska _ svenska _ engelska
Om du upplever att du blivit fel bemött inom hälsovården kan du ta kontakt med patientombudsmannen (potilasasiamies).
Arbetsgivaren arrangerar logi för merparten av arbetstagarna, och man strävar efter att ordna inkvartering så nära bygget som möjligt.
Läs noga anvisningarna om ansökning från den branschspecifika myndigheten.
Om den asylsökande beviljas uppehållstillstånd och är fast bosatt i Finland har han eller hon rätt till finskt socialskydd.
du äger minst 50 % av bostaden
InfoFinland är en mångsidig webbplats som sammanställer viktig information för personer som planerar att flytta till Finland eller som redan bor här.
Information om de samiska språkenfinska _ svenska
Mer information om äktenskapsförord får du på InfoFinlands sida Äktenskapsförord.
Arbets- och näringsbyrån eller TE-byrån (TE-toimisto) ger dig handledning i jobbsökningen och information om lediga jobb och tillgängliga utbildningar.
Handikappade personer har rätt att leva ett normalt liv, till exempel studera, arbeta och bilda familj.
För att få tillståndet krävs inga andra skäl, som till exempel arbete eller studier.
Säkerställ att du har följande när du kommer till Finland för att studera:
Förlängning av visum i Finlandfinska _ svenska _ engelska
Om du har frågor om den grundläggande utbildningen kan du kontakta skolbyrån.
Om du har kommit till Finland som kvotflykting och vill att finska staten bekostar resan för dina familjemedlemmar ska du ta kontakt med Röda Korsets beredskapsenhet som sätter igång researrangemangen.
Arbets- och näringsbyrån köper den yrkesinriktade arbetskraftsutbildningen av olika läroanstalter och företag.
skal från frukt och grönsaker
Du kan komma till Finland som utbytesstudent.
Om du vill skaffa dig praktiska kunskaper på en arbetsplats, är ett utbildningsavtal ett bra alternativ för ett läroavtal.
Köpcentret Grani
Svaret skickas till din e-post och publiceras på tjänstens webbplats.
Du kan även ansöka till utbildningen själv.
Ta också del av InfoFinlands sidor Ekonomiskt stöd till familjer och Vård av barnet.
Om det finns problem i familjen kan barnet själv be om vård utom hemmet.
På stadens webbplats finns skolornas kontaktuppgifter och mer information om anmälan.
Esbo handikappservice
Om du har symtom kan du utan remiss besöka Helsingfors poliklinik för könssjukdomar mån–fre kl. 8–12.
Esbo stads handikappservice
Handboken Jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
Barnskyddslagen gäller alla barn som bor i Finland oavsett deras nationalitet, religion eller kultur.
Tfn 09 276 62 899
Läs mer: Studier som hobby.
I dagvården lär barnet känna den finländska kulturen, lär sig det finska språket och verkar i en social grupp.
Lektionerna är vanligen 45 minuter långa.
Om du inte har hemvist i Finland eller något annat land inom EES, måste du registrera din företagsverksamhet i Patent- och registerstyrelsens handelsregister innan du ansöker om uppehållstillstånd för företagare.
Tjänsten har öppet måndag till fredag kl. 8–16.
Barn under 18 år ska alltid ha en minst en vårdnadshavare.
Stödets omfattning beror på den boendes behov.
Detta är dock det sista alternativet.
Om din maka/make har uppehållstillstånd i Finland på grund av internationellt skydd och flyktingstatus, kan du få uppehållstillstånd i Finland på grund av familjeband.
Gå och titta på bostaden innan du hyr den.
Föreningarfinska _ svenska
Lägg till bilagorna till ansökningen.
Detta innebär att modern ensam bestämmer om barnets angelägenheter även om föräldrarna bor tillsammans.
För praktik till Finland
Kristjänsterfinska _ svenska
I ansökningen ska du motivera varför du borde antas till utbildningen.
De presenterar konst, historia, natur, någon person eller ett specialområde.
du är själv fast bosatt i bostaden
Blanketterna finns på verksamhetsställena och på internet.
Information om konsumenträttigheterfinska _ svenska _ engelska
Läs mer: Yrkesutbildning
Om du drabbas av en akut krissituation, såsom att en närstående avlider eller på grund av familjevåld, kan du kontakta social- och krisjouren (sosiaali- ja kriisipäivystys).
Du kan även boka en telefontid vid FPA.
Du kan besöka en privat tandläkare även om du inte har rätt att anlita tjänster inom den offentliga hälso- och sjukvården.
Barnskyddet är baserat på lag
Tjänsterna är kostnadsfria.
Om du är studerande kan du söka en hyresbostad som är avsedd särskild för studerande. Studentbostäderna har oftast en lägre hyra än andra bostäder.
Om du är EU-medborgare och flyttar till Finland för att bo hos en familjemedlem ska du ansöka om registrering av uppehållsrätten för EU-medborgare på grund av familjeband i tjänsten Enter Finland eller på Migrationsverkets (Maahanmuuttovirasto) tjänsteställe.
En del människor, till exempel åldringar och handikappade, har svårt att klara av de dagliga sysslorna utan hjälp.
Små barn kan delta i verksamheten tillsammans med sin förälder eller vårdare.
Du kan kontakta intressanta organisationer direkt och fråga om de har lediga jobb.
Information om sjukförsäkringfinska _ svenska _ engelska
Flyktingrådgivningen
Orsaker till förföljelse kan vara etniskt ursprung, religion, medborgarskap, tillhörighet till en viss grupp i samhället eller politiska åsikter.
Telefon: 0295 025 500
Boka en tid vid Migrationsverkets tjänsteställe på Migrationsverkets webbplats.
Företagshälsovård kan ordnas på den lokala hälsovårdscentralen (terveyskeskus) eller till exempel en privat läkarstation.
linkkiFinlands översättar- och tolkförbund:
Du hittar mer information om religionsutövning i Finland på InfoFinlands sida Kulturer och religioner i Finland.
Ordlista om boendefinska
Mer information om detta hittar du på InfoFinlands sida Kan jag förlora mitt uppehållstillstånd?.
Esbo moderna konstmuseum EMMA är ett av Finlands största konstmuseer.
Huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors.
Du kan emellertid behöva en standardblankett som används som översättningsstöd som bilaga till en allmän handling.
Det består av fem dokument som har till syfte att hjälpa arbetstagare och studerande att presentera sitt kunnande i Europa.
Många museer ger rabatt på inträdesavgiften till vissa grupper.
Du måste då betala mäklararvode till mäklaren.
Till exempel uppmuntras unga vuxna att bli självständiga och flytta hemifrån.
Vanligen kan du arbeta högst 25 timmar i veckan.
grundläggande service, rättsskydd och tillstånd
Vid behov skriver tandläkaren en remiss till specialtandvården.
Registrering av utlänningar på skattebyrånfinska _ svenska _ engelska
Fackförbund
Mer information om uppehållstillstånd för studerande och om den sjukförsäkring som krävs för att få uppehållstillstånd får du på InfoFinlands sida Att studera i Finland eller på Migrationsverkets (Maahanmuuttovirasto) webbplats.
Barn och ungdomar kan studera musik vid Grankulla musikinstitut och bildkonst vid Grankulla konstskola.
Feedback till stadens ämbetsverk och inrättningarfinska _ svenska _ engelska
För detta behöver du barnets födelseattest från magistraten.
boende
Du får mer information om att ansöka om fortsatt uppehållstillstånd på InfoFinlands sida Fortsatt uppehållstillstånd.
Information om beslutet ges genom tolkning eller översättning.
Andra universitetsstudier leder inte till ett visst yrke.
Tillstånd för företagare som är bosatta utanför EES-områdetfinska _ svenska _ engelska
Tillstånd eller anmälan
Om du vill kan du efter magisterexamen söka till fortsatta studier.
I Karleby finns mångsidiga motionsmöjligheter året runt.
Lapplands TE-byrå betjänar kunderna per telefon måndagar, onsdagar, och torsdagar kl. 8–16.15 samt tisdagar och fredagar kl. 9–16.15 på numret 0295 039 501
avläggande av delar av ovan nämnda examina.
I Finland utförs egentliga elarbeten endast av personer som är yrkesutbildade inom elbranschen.
Om du är medborgare i något nordiskt land behöver du inte uppehållstillstånd i Finland.
Hur söker du dig till rehabilitering
I Finland dricker också vuxna ofta mjölk.
Läs mer: Fritidsverksamhet för barn och unga.
Mer information om reglerna i Finland ges av Livsmedelssäkerhetsverket Evira.
I Helsingfors finns ett stort antal olika föreningar, till exempel kulturföreningar och idrottsorganisationer.
Du hittar kontaktuppgifterna på webbplatsen ihmiskauppa.fi.
Juridisk hjälp kan du be om vid rättshjälpsbyrån (oikeusaputoimisto).
Servicepunkt för socialarbete och socialhandledningfinska _ svenska _ engelska
Napapiirin Residuum
Det lönar sig att söka till vissa utbildningar på främmande språk i den gemensamma ansökan i januari.
Vid behov får du rådgivning om hur du ansöker om utkomststödet hos FPA, socialbyrån i din hemkommun eller en rådgivning för invandrare.
Erkännande av examen
Om fadern inte erkänner sitt faderskap kan modern väcka talan för fastställande av faderskapet.
Brottsofferjouren
Du hittar kontaktuppgifterna till dem till exempel på Finlands översättar- och tolkförbunds webbplats.
Beroende på årstiden och området finns det olika aktivitetsmöjligheter.
Språkvalet kan påverka barnets möjligheter att studera olika språk i skolan.
Finska som andra språk i den grundläggande undervisningenfinska _ svenska
Programguideengelska
Beskattning
de inkomster som du har haft från början av året
I Finland ska man alltid på förhand komma överens om besök hos andra, även hos goda vänner.
I södra Finland reser man ibland också midsommarstången.
Socialbyråerna betjänar kommuninvånarna till exempel i följande ärenden:
Medling kan ofta vara nyttig och hjälpa er att komma överens i olika frågor utan rättegång.
De har tagit lån eller finansierat sin bostad på andra sätt.
mån–fre kl. 8.15–16.00
Många flygbolag erbjuder flyg från Finland till utlandet.
Bevis för yrkeskunnighet med fristående examen
Väestöliittos mentorskap i fråga om arbetskarriär är avsett för utbildade invandrare.
Din flytt till Finland kan betraktas som stadigvarande i följande situationer:
Åldringar kan använda tjänsterna vid de vanliga hälsostationerna.
Också myndigheterna måste följa lagen.
Områdeskoordinatorerfinska
Möjligheter att studera finska eller svenska
När du tar hand om en gammal eller sjuk anhörig eller en anhörig med funktionsnedsättning för att han eller hon ska kunna bo kvar i sitt hem, kan du ha rätt till stöd för närståendevård.
Om din bostad har skadats, till exempel till följd av brand eller vattenskada, kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna.
Huruvida du behöver ett uppehållstillstånd beror på i vilket land du är medborgare, varför du kommer till Finland och hur länge du ska stanna.
Be om kontaktuppgifterna till patientombudsmannen vid den vårdenhet där du har varit klient.
Skattebeloppet justeras i efterskott utgående från hur stora dina inkomster och avdrag verkligen har varit.
Allmän information om studier i finska och svenska i Finland hittar du på InfoFinlands sida Finska och svenska språket.
Mer information om medling i familjefrågor hittar du på InfoFinlands sida Skilsmässa.
I krigen förlorade Finland områden till Sovjetunionen.
När du är utomlands kan din sociala trygghet påverkas till exempel av att du inleder studier eller börjar arbeta.
Om du är företagare kan du bli medlem i företagarnas intressebevakningsorganisation Grankulla företagare rf som erbjuder sina medlemmar utbildning, nätverk och rådgivning.
Olika lån har olika villkor.
På webbtjänsten kan du söka och reservera material.
Magistraten utreder om du kan få en hemkommun registrerad.
Till dagvårdsplatser för verksamhetsåret som börjar i augusti ansöker man senast i slutet av mars.
Handikappade barns fritid
Barnet har rätt att få undervisning i sin egen religion i skolan.
Arbetspensionen intjänas med det egna lönearbetet och företagandet.
I Finland finns en lag om likabehandling, som föreskriver att arbetsgivaren ska övervaka att jämställdheten på arbetsplatsen realiseras och att ingen diskrimineras på arbetsplatsen.
Tfn 045 639 6274
Sexuell hälsa hos kvinnor
Du kan kontakta rådgivningen via den centraliserade telefontjänsten (06) 826 4477.
Makarna kan vara partiellt vårdlediga samtidigt så att den ena förkortar sin arbetstid från morgonen och den andra från eftermiddagen.
Utöver pension kan FPA betala ut bostadsbidrag till pensionstagare med låga inkomster.
På InfoFinlands sida Ansökan till utbildning finns information om hur du ansöker till utbildning på andra stadiet och högskoleutbildning i Finland.
Läs mer på InfoFinlands sida Stöd för vård av barn i hemmet.
Räntestöd beviljas för unga som skaffar sin första ägarbostad.
Om du har betalat för lite i skatt, blir du tvungen att betala kvarskatt (jäännösvero).
Förskoleundervisningen börjar i augusti och anmälan ska göras i februari.
Information om kontaktuppgifter finns på Vanda stads webbplats.
I Finland är nätspänningen 230 volt.
MoniNet är ett mångkulturellt center i Rovaniemi, Lappland. Det upprätthålls av föreningen Rovalan Setlementti ry.
Studerande
Vårdnadshavare till en finsk medborgarefinska _ svenska _ engelska
Ansökan till en yrkesinriktad vuxenutbildning
Information om tolktjänsterfinska
Mångsidiga övningar i finska språketfinska
Grankulla stad erbjuder olika tjänster för handikappade, till exempel hjälpmedel och dagverksamhet.
Läkaren skriver en remiss till det sjukhus där aborten görs.
Om du behöver psykisk hjälp och psykiskt stöd kan du kontakta hälsostationen.
fysiska symptom, utan att medicinska orsaker hittas för dessa
I en del kommuner kan du delta i integrationsutbildning på svenska.
Om du och din sambo är bosatta i olika stater anses gemensamt boende till exempel under semesterresor inte som en tillräcklig grund för beviljande av uppehållstillstånd.
Inkomsterna för din partner som är bosatt i Finland beaktas inte.
Badhuset/+simhallen Vesihiisifinska
Om du behöver rättshjälp, kan du kontakta Helsingfors rättshjälpsbyrå (Helsingin oikeusaputoimisto).
Medlingen är kostnadsfri.
Denna gräns mellan religionerna finns fortfarande, men med reformationen byttes den katolska tron till den lutherska.
Kommunerna är skyldiga att ordna många olika tjänster för sina invånare.
Var får jag hjälp?
Vuxengymnasiumfinska
Stöd och hjälp för handikappade invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ persiska _ arabiska _ kurdiska
Kommunerna måste tillhandahålla handikappade de tjänster som de behöver.
Privata servicehusfinska
När föräldrarna har kommit överens om barnets boende, vårdnad, umgängesrätt och underhållsbidrag kan socialväsendet på orten bekräfta avtalet.
Studieutbudet är väldigt mångsidigt.
Om bostaden har centralvärme, ingår uppvärmningen i allmänhet i hyran.
Vid rådgivningen följs moderns, fostrets och hela familjens hälsotillstånd under graviditeten.
I anslutning till TE-byrån finns ett rum där man kan uträtta ärenden på egen hand.
I Grankulla finns också privata tandläkare.
Din grundutbildning avgör till hurudan yrkesutbildning du kan söka och på vilket sätt ansökan sker.
I Helsingfors, Åbo, Tammerfors och Esbo får barn och gravida kvinnor samma hälso- och sjukvårdstjänster som övriga invånare.
Ekonomiskt stöd under den yrkesinriktade arbetskraftsutbildningen
Till exempel finns det information om kurserna i finska språket i Helsingfors, Tammerfors och Åbo i tjänsten Finnishcourses.fi.
Sexuell hälsa hos män
I Esbo finns flera bibliotek på olika håll i staden.
Preventivmedel säljs på apoteket.
Hur kan man minska mängden avfall?
Anmäl dig som arbetssökande i TE-byråns webbtjänst.
Om ett barn blir sjukt och behöver snabbt vård, ta kontakt med hälsostationen (terveysasema).
Många medborgarorganisationer och föreningar har särskilda ungdomsavdelningar som ordnar verksamhet för unga.
Information för flyktingarfinska _ engelska _ franska _ persiska _ arabiska _ kurdiska
Du kan ofta boka läkartiden via mödrarådgivningen.
Självrisktiden är vanligen den dag då du insjuknade och därpå följande nio vardagar.
Finland blev självständigt 1917.
linkkiArbets- och näringsministeriet:
Följ informationen på arbetsplatsen.
Om detta inte hjälper, kan du kontakta disponenten eller hyresvärden.
Serviceguide för handikappade invandrare(pdf, 797,26)finska _ engelska _ ryska _ arabiska
De sköter begravningsarrangemangen, som till exempel transporten av den avlidne.
Stödet är avsett för dem som har en hemkommun i Finland.
Finland har 5,5 miljoner invånare.
Konflikter med grannarna
Den är avsedd för de elever som ännu inte har särskilt bra kunskaper i finska.
linkkiAvfallsverksföreningen:
Om du vistas utomlands tillfälligt, det vill säga under ett år, betalar FPA vanligtvis din pension som vanligt.
Att studera i Finland
Hyresvärden har rätt att häva hyresavtalet om du inte betalar din hyra.
Att tvinga någon till äktenskap är ett brott i Finland.
Hälsostationernafinska _ svenska _ engelska
Hälsostationerna har öppet från måndag till fredag, vanligen kl. 8–16.
Kontaktuppgifter till enheten som väljer hyresgästerna, telefontid kl. 12–15:
Om till exempel utbildning i läs- och skrivkunnighet eller någon annan språkutbildning har godkänts till din integrationsplan, tas det inte ut någon avgift för studierna.
Du kan vända dig till diskrimineringsombudsmannen till exempel om du själv har råkat ut för etnisk diskriminering eller observerat att en annan person diskrimineras.
Fråga din arbetsgivare som hen använder tjänsten Enter Finland för arbetsgivare.
linkkiFaro:
Om din finländska arbetsgivare har sänt dig utomlands för att arbeta förlorar du inte ditt uppehållstillstånd i Finland även om du vistas utomlands på grund av arbetet i över två år.
Uleåborg
Dessutom övervakar riksdagen regeringens verksamhet.
Om familjen har barn under 18 år och äktenskapet slutar ska föräldrarna i samband med skilsmässan komma överens om följande:
Grankulla socialbyrå
Vinterkriget och fortsättningskriget
skattebyrån, om du behöver personbeteckningen för beskattningen.
Skattebyrån (verotoimisto) har ett serviceställe i centrala Helsingfors.
Ansökan kan även göras senare, men då tillämpas kravet på tillräcklig inkomst.
Vanligtvis kan man få FPA:s bidrag då de övriga inkomsterna är låga.
Detta får inte orsaka extra kostnader för patienten.
När du ansöker om ditt första uppehållstillstånd i Finland kan du även be om att bli registrerad i Finlands befolkningsdatasystem.
Om du har ett uppehållstillstånd för arbetstagare som endast gäller arbete för en viss arbetsgivare och du förlorar din arbetsplats, ska du ansöka om ett nytt uppehållstillstånd för arbetstagare eller ett uppehållstillstånd på andra grunder.
För att få bostadsbidrag måste du också du omfattas av den sociala tryggheten i Finland.
I vissa fall kan du alltså inte få webbankkoder även om du har ett bankkonto.
Anvisningar för jobbintervjunfinska _ svenska _ engelska
Du kan ansöka om finskt medborgarskap när du har fyllt 18 år, har bott permanent i Finland i tillräckligt många år, har nöjaktiga muntliga och skriftliga kunskaper i finska eller svenska eller motsvarande kunskaper i finskt eller finlandssvenskt teckenspråk och din identitet är tillförlitligt utredd.
Om du inte avbokar debiteras du på en avgift om 27 euro.
Barn
12–17 år och adoptivbarn till en finsk medborgare
Rehabilitering för gravt handikappade
Grunderna för antagning av studeranden beror på utbildningen.
Familjerådgivningfinska _ engelska
I Finland finns många patientföreningar som tillhandahåller information och rådgivning för människor med en viss sjukdom.
Samtal till Nollalinja är kostnadsfria och de syns inte i telefonräkningen.
Sådana stipendier är till exempel de som beviljats av staten, läroanstalter eller organisationer.
Också tillräckliga medel är en grund.
Föräldrapenning
Stadin aikuisopisto ordnar i vissa lekparker och familjehus kurser i finska för invandrarföräldrar.
Invandrartjänster
du har ett gemensamt barn med din sambo (då uteblir kravet på gemensamt boende under två års tid) eller
Om det finns minst tio anställda på en arbetsplats väljer dessa ut en arbetarskyddsfullmäktig som representerar dem.
Vid behov skriver läkaren en remiss till den psykiatriska polikliniken för dig.
Du kan även ansöka till yrkesutbildning för vuxna.
Läs mer på InfoFinlands sida Gymnasieförberedande utbildning.
Val av vigselform
Övernattningsalternativ i Karlebyfinska _ svenska _ engelska
Modersmålsprovet är ett obligatoriskt prov i studentexamen.
Privata hyresbostäder
En familjebostad är en omöblerad lägenhet som endast hyrs ut till personer i samma hushåll.
Du kan grunda ett aktiebolag antingen själv eller tillsammans med andra delägare.
Förmodligen får du en tid snabbare på en privat hälsostation än inom den offentliga hälsovården.
Du kan också boka tid hos en privat tandläkare.
Stödet kommer från samhället i form av den sociala tryggheten.
Kom ihåg att kontrollera också det nya beskattningsbeslutet.
Du kan utarbeta en integrationsplan t.ex. med en arbetskraftsrådgivare vid arbets- och näringsbyrån, alltså TE-byrån (TE-toimisto), eller med en socialarbetare på socialbyrån.
Du har rätt att utnyttja de offentliga hälsovårdstjänsterna om du har hemkommun i Finland.
Mer information om dessa språk får du på webbplatsen för Forskningscentralen för de inhemska språken.
Det är lättare att söka jobb om du vet hur en examen som du avlagt utomlands motsvarar en finländsk examen.
På InfoFinlands sida Utbildning i Grankulla finns information om dagvård för barn.
I Finland ägs cirka 70 procent av idrottsanläggningarna av kommunerna.
Jag är lärare / ingenjör / studerande.
Äktenskapsförord är frivilligt.
Även om finländarna i allmänhet behärskar engelska relativt väl har du ändå mycket nytta av att kunna finska eller svenska.
Telefon: 040 806 8101
Om du inte kan betala dina räkningar eller skulder då de förfaller, ska du kontakta skuldrådgivningen (velkaneuvonta).
Du kan söka svenskspråkiga högskoleutbildningar via tjänsten Opintopolku.fi.
Information om småbarnspedagogikfinska _ svenska _ engelska
Köp endast sådana saker du behöver.
Motionsrekommendationerfinska _ engelska
Om du vill förbättra dina kunskaper i finska eller svenska innan du söker till ett gymnasium, kan du söka till en förberedande gymnasieutbildning.
Hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
Studentbostäderna är oftast billigare än bostäderna på den öppna marknaden.
Boka en tid på mödrarådgivningen.
Grunddagpenningfinska _ svenska _ engelska
Anmäl dig till husets ägare.
En läkare eller någon annan yrkesutbildad person avgör detta.
Om du behöver stöd för din integration, utarbetas en integrationsplan för dig efter den inledande kartläggningen.
Observera att officiella handlingar som tagits med från utlandet ska vara legaliserade och i original samt översatta till finska, svenska eller engelska.
faderskapspenning.
Privat tandvård är dyrare än offentlig tandvård.
Handikappades rättigheter
Enligt Finlands lag är äktenskapet (avioliitto) ett lagstadgat förhållande mellan två människor.
På gymnasiet kan man även höja vitsorden i sitt avgångsbetyg eller studera enskilda ämnen.
Om barnet inte kan få krävande medicinska rehabilitering från FPA, ska rehabiliteringen ordnas av hemkommunen.
att slå, sparka och knuffa
linkkiBortförda barn rf:
Det självständiga Finland blev en republik där lagarna stiftas av en folkvald riksdag.
Du kan även studera språket på Internet.
Hälsovårdstjänster ges i Finland på finska och svenska.
Om du inte har en finländsk personbeteckning, är ditt bibliotekskort i kraft ett år i taget.
Tänk på att frivilligarbete kan påverka din arbetslöshetsförsäkring.
Påsen tillsluts noga.
Olika läkarstationer erbjuder olika tjänster.
Förnamnen ska vara förenliga med Finlands namnlag.
Information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb?
Svenskspråkiga yrkesläroanstalter och gymnasieskolor finns i svenskspråkiga och tvåspråkiga kommuner och i en del finskspråkiga kommuner.
Uppsägningstiden är den tid som arbetstagaren är skyldig att arbeta innan arbetet upphör.
Boendetjänster för handikappadefinska _ svenska _ engelska
Finland ligger i Nordeuropa.
Under Ryssland blev Finland ett speciellt område som utvecklades på kejsarens order.
Om du vill ta en personförsäkring i ett finländskt försäkringsbolag ska du vanligtvis ha ett finländskt FPA-kort.
Ibland krävs att du lyckas tillräckligt bra med dina studier för att du ska få ett stipendium.
Underhållsbidraget har på grund av förälderns ekonomiska situation fastställts till ett belopp som underskrider underhållsstödet.
Uppehållstillstånd för studerande från andra EU-länder
Yrkeshögskoleexamen kan avläggas på 3,5–4,5 år.
Helsingfors är även ett viktigt centrum för affärs- och kulturlivet.
Gymnasiet ger förberedande utbildning till exempel för yrkeshögskola och universitet.
en talskada
Om originalspråket för ditt betyg inte är finska, svenska eller engelska behöver du vanligtvis en officiell översättning av handlingarna som görs av en auktoriserad översättare.
Vem som helst kan studera vid dessa.
Information om tjänster för äldrefinska _ svenska _ engelska
Det är bra att förvara filten till exempel i närheten av spisen.
Inom företagshälsovården har arbetstagaren tillgång till hälsovårdarens, företagsläkarens och företagspsykologens tjänster.
Om du flyttar utomlands
Att låna material
Om du eller din familj har utgifter på grund av särskilda behov, för vilka du inte kan få grundläggande utkomststöd, kan socialbyrån i din hemkommun bevilja kompletterande och förebyggande utkomststöd (täydentävä ja ehkäisevä toimeentulotuki).
Tfn 050 300 6093
Om du kommer till Finland för att studera kan du få en studentbostad där du får bo så länge som dina studier i Finland pågår.
Förskoleundervisningen ordnas av kommunerna och är kostnadsfri för familjen.
Vård av barn
Du kan rösta i kommunalvalet om:
Information om diskrimineringfinska _ svenska _ engelska
Hedersrelaterat våld
Att bo i en bostadsrättsbostad är ett alternativ till att köpa eller hyra sin bostad.
På beskattningen inverkar också huruvida din arbetsgivare är ett finländskt eller ett utländskt företag.
Det är lättast om operationen görs innan graviditeten har börjat, men den kan också göras i mitten av graviditeten.
Om du bor i östra Helsingfors, sydöstra Helsingfors, nordöstra Helsingfors eller norra Helsingfors hittar du hälsovårdscentraljouren vid Malms sjukhus.
Besläktade språk är till exempel estniska och ungerska.
Besöksadress:
Fennovoima bygger kärnkraftverksenheten Hanhikivi 1 i Pyhäjoki.
Helsingfors stad hjälper arbetslösa helsingforsare att hitta jobb eller utbildning.
vid social delaktighet,
Du kan byta ut ditt körkort till ett finskt körkort på Ajovarmas serviceställe.
Barnet kan också få hjälpmedel om han eller hon inte kan studera utan dem eller om det är mycket svårt utan dem.
att bevittna våldsamma situationer
om du redan har fött fyra barn
Stödet består antingen av pengar eller tjänster.
Vinter
Lönen kan innehålla olika förmåner.
du är medborgare i ett nordiskt land
Om du misstänker att du har en könssjukdom kan du boka en läkartid på hälsostationen eller en privat läkarstation.
Finskans uttal är mycket regelbundet.
Sådana är till exempel många idrotts- och simhallar och andra idrottsanläggningar, såsom fotbollsplaner och skridskobanor.
Du kan själv välja om du vill ta ut 25 procent eller 50 procent av beloppet på din månatliga arbetspension.
Om du behöver mer information om legalisering av handlingar, kontakta magistraten eller utrikesministeriet i ditt eget land.
För att få en inledande kartläggning gjord, ska du anmäla dig som arbetssökande via Internet på adressen te-palvelut.fi.
Prepaid-kortet är i förväg laddat med en summa som man sedan kan ringa för.
Dessa uppgifter är bland annat namn, födelsedatum, medborgarskap, kön och adress.
Fler än 400 000 finländare lämnade de förlorade områdena och kom som flyktingar till övriga delar av landet.
I Kelviå, ca 10 km norrut från Karleby, finns Toivonen djurpark och drängmuseum.
Anmäl diskrimineringfinska _ svenska _ engelska
Verksamheten i öppna daghem och invånarparker är kostnadsfri och du behöver inte anmäla dig på förhand.
Du kan ändå behöva ett visum.
Läs mera om privatvårdsstöd på Fpa:s sidor.
Andra religiösa samfund i Finland är till exempel Katolska kyrkan i Finland, Pingstkyrkan i Finland, Frikyrkan i Finland, Adventkyrkan i Finland, mormonkyrkan och Jehovas vittnen.
IHH – serviceställe för dig som flyttar till Finland engelska
Du ska vanligtvis även kunna visa ditt betalningsbeteende, dvs. uppgifter som visar att du har betalat dina räkningar och inte har några betalningsanmärkningar.
Det är tillåtet att spela in material på offentliga platser, för inspelning i privata lokaler ska tillstånd inhämtas.
Föreningens styrelse
Borgmästaren och stadens aktörer ordnar boendemöten runtom i Helsingfors för invånarna där man berättar om och diskuterar stadens ärenden.
Vem som helst kan studera vid en öppen högskola.
Förvara hyresavtalet noga.
Öppna linjen: 09 7562 2260
Hjälp för unga
