gör ansökan inom tre månader efter datumet för inresa .
en del tolkcentraler har jour på veckoslut samt kvällar och nätter .
kan den ena sambon inte få änkepension om den andra sambon dör .
fundera också på om du har tillräckliga yrkeskunskaper och erfarenhet .
Karleby verksamhetsställe
transporttjänster
använd inte elapparater som är i dåligt skick eller vars sladd är trasig .
Nuortenkatu 11
läs mer på InfoFinlands sida Tjänster för handikappade .
om du kommer som flykting till Finland ska du komma överens om en hälsokontroll med utlänningsbyrån .
Ansvarsområdena för arbetarskydd ger både arbetstagare och arbetsgivare råd i frågor som gäller arbetets säkerhet och hälsa samt i frågor som rör anställningsvillkor .
är fadern förpliktad att delta i underhåll av barnet
kvotflyktingar
faderskapsledighet
handläggning av ansökan om registrering av uppehållsrätt är avgiftsbelagd .
har det uppehållstillstånd ( oleskelulupa ) som krävs och
_ holländska _ kroatiska _ rumänska _ ungerska _ japanska _ italienska
myndigheter som utfärdar Apostilleintyg finns i alla länder som är anslutna till Haagkonventionen .
barnen har ofta en och samma lärare under de sex första skolåren .
FPA:s kunder är alla personer som bor i Finland och utomlands och som omfattas av socialskyddet i Finland .
om det till exempel anges i hyresavtalet att det är förbjudet att röka i bostaden , kan du inte röka i ditt hem .
om äktenskapet till exempel har varat under fem år delas egendomen inte nödvändigtvis jämnt .
Barnbidraget för det första barnet uppgår till cirka 100 euro per månad .
Jorvs sjukhus
i Finland visas filmerna oftast på originalspråket .
arbets- och näringsbyråerna och kommunerna tillhandahåller invandrarrådgivning .
behovsprövad rehabiliteringfinska _ svenska
om du inte tar emot platsen i tid , förlorar du den .
när du inleder företagsverksamheten har du många skyldigheter , bland annat ska du registrera företaget och ordna beskattning och bokföring .
om du redan är i Finland och får ett negativt beslut om uppehållstillstånd från Migrationsverket ( Maahanmuuttovirasto ) , måste du antingen lämna Finland eller överklaga beslutet .
till ansökan om uppehållstillstånd för arbetstagare ska du bifoga blanketten TEM054 som din arbetsgivare fyller i och undertecknar .
till exempel på Helsingfors stads webbplats finns en färdig blankett , ett responssystem ( palautejärjestelmä ) .
om din bostad har skadats till exempel till följd av brand eller vattenskada kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna .
när ni kräver bodelning förordnar tingsrätten en bodelningsman som delar egendomen .
Sanduddsgatan 5 B
du hittar kontaktuppgifterna på Sopu @-@ arbetets webbplats .
arbetstagare , företagare , studerande , flykting , asylsökande eller en familjemedlem till en person bosatt i Finland hittar information speciellt om sin egen situation på dessa sidor i Infobanken .
du får hjälp med spelproblem vid A @-@ kliniker ( A @-@ klinikka ) , mentalvårdsbyråer ( mielenterveystoimisto ) och hälsovårdscentralen ( terveyskeskus ) .
om du blir bostadslös , kontakta Esbo stads verksamhetsställe för vuxensocialarbete .
tjänsterna och priserna i olika flyttfirmor kan variera stort och därför lönar det sig att jämföra .
i Vanda finns 10 bibliotek ( kirjasto ) och två bokbussar ( kirjastoauto ) .
Infomötena är avgiftsfria .
det kan vara fördelaktigt att kunna svenska när du söker jobb .
startpenning
ensamboende eller
stöd för skolresor
i Finland kan du avbryta en graviditet i tidigt skede i följande fall :
om dina studier fortsätter men uppehållstillståndet håller på att gå ut ska du ansöka om fortsatt uppehållstillstånd .
information om priser på sålda bostäderfinska _ svenska
Mun- och tandhälsovårdenfinska _ svenska _ engelska
linkkiHelsingforsregionens miljötjänster :
när din examensnivå har jämställts med en finländsk högskoleexamen , kan du söka till uppgifter som kräver den nivå på högskoleexamen som du har .
Skriv alltid ett skriftligt anställningsavtal innan du börjar på ett nytt jobb .
i de allra nordligaste delarna av Finland går solen inte alls ner i början av sommaren .
någon hotar dig eller din familj med våld
information om boendefinska _ engelska
barnen äter en varm måltid i skolan .
mer information om juristtjänster och rättshjälp hittar du på InfoFinlands sida Behöver du en jurist ? .
Heminkvarteringengelska _ franska _ spanska _ kinesiska _ tyska _ portugisiska _ italienska
när du ansöker om startpeng undersöker TE @-@ byrån om företagandet är ett lämpligt alternativ för dig .
finländare väntar vanligtvis att samtalspartnern har sagt sitt innan de själva tar till ordet .
linkkiFörbundet för Steinerpedagogik :
om du inte förstår finska eller det finska teckenspråket kan du också behöva en annan tolk .
du kan söka olika föreningar i patent- och registerstyrelsens tjänst Föreningsregistret .
i arbetsavtalet fastställs arbetsuppgifterna och lönen samt andra förmåner och villkor .
om din arbetserfarenhet i Finland är kort eller om din finska ännu inte är så bra , kan frivilligarbete vara ett bra sätt att få fotfäste i arbetslivet och förbättra språkkunskaperna .
boende i bostadsrättsbostad
( det är bra att veta att stadigvarande boende definieras på olika sätt i olika lagar .
under prövotiden kan arbetstagaren och arbetsgivaren häva arbetsavtalet utan uppsägningstid .
tfn 045.134.1711
Prästgårdsgränden 5
läroplikten upphör när barnet har fullgjort hela lärokursen för den grundläggande utbildningen eller det har förflutit tio år sedan läroplikten började .
företagare måste inte ordna företagshälsovård för sig själv , men däremot måste de ordna det för sina anställda .
om du vill att en mäklare söker en lämplig hyresbostad åt dig , ska du ingå ett skriftligt uppdragsavtal ( toimeksiantosopimus ) med mäklaren .
Guide om att grunda ett företagfinska _ engelska _ kinesiska
linkkiEvangelisk @-@ lutherska kyrkan i Finland :
bostadslån
om du upprepade gånger bryter mot husets ordningsregler har hyresvärden rätt att häva hyresavtalet .
den som är en enskild näringsidkare beskattas på så sätt att alla inkomster som återstår efter att man har dragit av kostnaderna för företagsverksamheten är beskattningsbara inkomster .
Tillstånet kan dras tillbaka om du permanent flyttar från Finland , uppehåller dig utomlands kontinuerligt i minst två år eller har lämnar felaktiga uppgifter då du ansökt om tillståndet .
detta är det bra att beakta när du väljer företagsform .
gravplats
de flesta jobben är dolda jobb .
för vilka studier kan man få arbetslöshetsförmån ?
kontrollera detta med din arbetsgivare .
Nattcentret Kalkkersfinska
både offret och förövaren kan få hjälp .
finska medborgare kan i Finland dömas för brott som begåtts utomlands .
till exempel utbytesstuderande får inte finskt studiestöd .
du ska också ha en giltig trafikförsäkring ( liikennevakuutus ) för din bil i Finland .
vardera maken ansvarar ensam för den skuld som de har tagit före äktenskapet eller under det .
Finlands historia är en berättelse om handelsvägar , möten mellan kulturer och livet intill stora grannar .
undervisning i den egna religionenfinska
brådskande psykiatrisk sjukvård ges på jourenheter vid psykiatriska sjukhus .
Företagsfinland
tfn ( 09 ) 622.4322
stöd och handledning för ungafinska _ engelska
Flerspråkiga biblioteket
närskolan är oftast den skola som ligger närmast barnets hem .
du kan också köpa avgiftsbelagda kanaler .
du måste ha med ett ID @-@ kort när du röstar .
fråga mer på din hälsostation .
om du vistas i Finland i mer än sex månader , ska du i allmänhet betala skatt på din lön till Finland .
när du ansöker om startpenning utreder arbets- och näringsbyrån om företagande är ett lämpligt alternativ för dig .
för att kunna ansöka om en hyresbostad hos staden , måste du ha uppehållstillstånd för minst ett år .
information om kurser i skidåkning , om att hyra skidor och om skidspår finns till exempel på Suomen Latu ry:s webbplats på finska .
förberedande utbildning inför yrkesutbildning
Finest sänder radioprogram på estniska .
experterna där hjälper dig att utveckla affärsidén . du får hjälp med att utarbeta preliminära marknadsundersökningar , lönsamhetskalkyler och en kartläggning om tillgången till finansiering .
olika instanser anordnar företagarkurser och informationsmöten som man har mycket nytta av om man vill starta ett företag .
begäran om prövning kan ställas på vilken magistrat som helst .
tfn 016.3222.570 .
du ska ta pillret så snart som möjligt efter samlaget , i regel senast inom 72 timmar .
Karlebygatan 74
Dagvårdsavgifterfinska _ svenska _ engelska
om du upplever att du blivit fel bemött inom hälsovården kan du ta kontakt med patientombudsmannen ( potilasasiamies ) .
arbetsgivaren arrangerar logi för merparten av arbetstagarna , och man strävar efter att ordna inkvartering så nära bygget som möjligt .
läs noga anvisningarna om ansökning från den branschspecifika myndigheten .
om den asylsökande beviljas uppehållstillstånd och är fast bosatt i Finland har han eller hon rätt till finskt socialskydd .
du äger minst 50 % av bostaden
InfoFinland är en mångsidig webbplats som sammanställer viktig information för personer som planerar att flytta till Finland eller som redan bor här .
information om de samiska språkenfinska _ svenska
mer information om äktenskapsförord får du på InfoFinlands sida Äktenskapsförord .
arbets- och näringsbyrån eller TE @-@ byrån ( TE @-@ toimisto ) ger dig handledning i jobbsökningen och information om lediga jobb och tillgängliga utbildningar .
handikappade personer har rätt att leva ett normalt liv , till exempel studera , arbeta och bilda familj .
för att få tillståndet krävs inga andra skäl , som till exempel arbete eller studier .
Säkerställ att du har följande när du kommer till Finland för att studera :
förlängning av visum i Finlandfinska _ svenska _ engelska
om du har frågor om den grundläggande utbildningen kan du kontakta skolbyrån .
om du har kommit till Finland som kvotflykting och vill att finska staten bekostar resan för dina familjemedlemmar ska du ta kontakt med Röda Korsets beredskapsenhet som sätter igång researrangemangen .
arbets- och näringsbyrån köper den yrkesinriktade arbetskraftsutbildningen av olika läroanstalter och företag .
skal från frukt och grönsaker
du kan komma till Finland som utbytesstudent .
om du vill skaffa dig praktiska kunskaper på en arbetsplats , är ett utbildningsavtal ett bra alternativ för ett läroavtal .
Köpcentret Grani
Svaret skickas till din e @-@ post och publiceras på tjänstens webbplats .
du kan även ansöka till utbildningen själv .
ta också del av InfoFinlands sidor Ekonomiskt stöd till familjer och vård av barnet .
om det finns problem i familjen kan barnet själv be om vård utom hemmet .
på stadens webbplats finns skolornas kontaktuppgifter och mer information om anmälan .
Esbo handikappservice
om du har symtom kan du utan remiss besöka Helsingfors poliklinik för könssjukdomar mån @-@ fre kl . 8 @-@ 12 .
Esbo stads handikappservice
Handboken jobba i Finlandfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ kinesiska _ arabiska _ kurdiska _ tyska _ thai _ vietnamesiska
barnskyddslagen gäller alla barn som bor i Finland oavsett deras nationalitet , religion eller kultur .
tfn 09.276.62.899
läs mer : studier som hobby .
i dagvården lär barnet känna den finländska kulturen , lär sig det finska språket och verkar i en social grupp .
Lektionerna är vanligen 45 minuter långa .
om du inte har hemvist i Finland eller något annat land inom EES , måste du registrera din företagsverksamhet i Patent- och registerstyrelsens handelsregister innan du ansöker om uppehållstillstånd för företagare .
tjänsten har öppet måndag till fredag kl . 8 @-@ 16 .
barn under 18 år ska alltid ha en minst en vårdnadshavare .
Stödets omfattning beror på den boendes behov .
detta är dock det sista alternativet .
om din maka / make har uppehållstillstånd i Finland på grund av internationellt skydd och flyktingstatus , kan du få uppehållstillstånd i Finland på grund av familjeband .
gå och titta på bostaden innan du hyr den .
föreningarfinska _ svenska
lägg till bilagorna till ansökningen .
detta innebär att modern ensam bestämmer om barnets angelägenheter även om föräldrarna bor tillsammans .
för praktik till Finland
Kristjänsterfinska _ svenska
i ansökningen ska du motivera varför du borde antas till utbildningen .
de presenterar konst , historia , natur , någon person eller ett specialområde .
du är själv fast bosatt i bostaden
Blanketterna finns på verksamhetsställena och på internet .
information om konsumenträttigheterfinska _ svenska _ engelska
läs mer : yrkesutbildning
om du drabbas av en akut krissituation , såsom att en närstående avlider eller på grund av familjevåld , kan du kontakta social- och krisjouren ( sosiaali- ja kriisipäivystys ) .
du kan även boka en telefontid vid FPA .
du kan besöka en privat tandläkare även om du inte har rätt att anlita tjänster inom den offentliga hälso- och sjukvården .
barnskyddet är baserat på lag
tjänsterna är kostnadsfria .
om du är studerande kan du söka en hyresbostad som är avsedd särskild för studerande . Studentbostäderna har oftast en lägre hyra än andra bostäder .
om du är EU @-@ medborgare och flyttar till Finland för att bo hos en familjemedlem ska du ansöka om registrering av uppehållsrätten för EU @-@ medborgare på grund av familjeband i tjänsten Enter Finland eller på Migrationsverkets ( Maahanmuuttovirasto ) tjänsteställe .
en del människor , till exempel åldringar och handikappade , har svårt att klara av de dagliga sysslorna utan hjälp .
små barn kan delta i verksamheten tillsammans med sin förälder eller vårdare .
du kan kontakta intressanta organisationer direkt och fråga om de har lediga jobb .
information om sjukförsäkringfinska _ svenska _ engelska
Flyktingrådgivningen
orsaker till förföljelse kan vara etniskt ursprung , religion , medborgarskap , tillhörighet till en viss grupp i samhället eller politiska åsikter .
telefon : 0295.025.500
boka en tid vid Migrationsverkets tjänsteställe på Migrationsverkets webbplats .
företagshälsovård kan ordnas på den lokala hälsovårdscentralen ( terveyskeskus ) eller till exempel en privat läkarstation .
linkkiFinlands översättar- och tolkförbund :
du hittar mer information om religionsutövning i Finland på InfoFinlands sida kulturer och religioner i Finland .
Ordlista om boendefinska
mer information om detta hittar du på InfoFinlands sida Kan jag förlora mitt uppehållstillstånd ? .
Esbo moderna konstmuseum EMMA är ett av Finlands största konstmuseer .
huvudstadsregionens skattebyrå ligger på Alexandersgatan 9 i Gloet i Helsingfors .
du kan emellertid behöva en standardblankett som används som översättningsstöd som bilaga till en allmän handling .
det består av fem dokument som har till syfte att hjälpa arbetstagare och studerande att presentera sitt kunnande i Europa .
många museer ger rabatt på inträdesavgiften till vissa grupper .
du måste då betala mäklararvode till mäklaren .
till exempel uppmuntras unga vuxna att bli självständiga och flytta hemifrån .
vanligen kan du arbeta högst 25 timmar i veckan .
grundläggande service , rättsskydd och tillstånd
vid behov skriver tandläkaren en remiss till specialtandvården .
registrering av utlänningar på skattebyrånfinska _ svenska _ engelska
fackförbund
mer information om uppehållstillstånd för studerande och om den sjukförsäkring som krävs för att få uppehållstillstånd får du på InfoFinlands sida Att studera i Finland eller på Migrationsverkets ( Maahanmuuttovirasto ) webbplats .
barn och ungdomar kan studera musik vid Grankulla musikinstitut och bildkonst vid Grankulla konstskola .
Feedback till stadens ämbetsverk och inrättningarfinska _ svenska _ engelska
för detta behöver du barnets födelseattest från magistraten .
boende
du får mer information om att ansöka om fortsatt uppehållstillstånd på InfoFinlands sida Fortsatt uppehållstillstånd .
information om beslutet ges genom tolkning eller översättning .
andra universitetsstudier leder inte till ett visst yrke .
tillstånd för företagare som är bosatta utanför EES @-@ områdetfinska _ svenska _ engelska
tillstånd eller anmälan
om du vill kan du efter magisterexamen söka till fortsatta studier .
i Karleby finns mångsidiga motionsmöjligheter året runt .
Lapplands TE @-@ byrå betjänar kunderna per telefon måndagar , onsdagar , och torsdagar kl . 8 @-@ 16.15 samt tisdagar och fredagar kl . 9 @-@ 16.15 på numret 0295.039.501
avläggande av delar av ovan nämnda examina .
i Finland utförs egentliga elarbeten endast av personer som är yrkesutbildade inom elbranschen .
om du är medborgare i något nordiskt land behöver du inte uppehållstillstånd i Finland .
hur söker du dig till rehabilitering
i Finland dricker också vuxna ofta mjölk .
läs mer : fritidsverksamhet för barn och unga .
mer information om reglerna i Finland ges av Livsmedelssäkerhetsverket Evira .
i Helsingfors finns ett stort antal olika föreningar , till exempel kulturföreningar och idrottsorganisationer .
du hittar kontaktuppgifterna på webbplatsen ihmiskauppa.fi .
juridisk hjälp kan du be om vid rättshjälpsbyrån ( oikeusaputoimisto ) .
servicepunkt för socialarbete och socialhandledningfinska _ svenska _ engelska
Napapiirin Residuum
det lönar sig att söka till vissa utbildningar på främmande språk i den gemensamma ansökan i januari .
vid behov får du rådgivning om hur du ansöker om utkomststödet hos FPA , socialbyrån i din hemkommun eller en rådgivning för invandrare .
erkännande av examen
om fadern inte erkänner sitt faderskap kan modern väcka talan för fastställande av faderskapet .
Brottsofferjouren
du hittar kontaktuppgifterna till dem till exempel på Finlands översättar- och tolkförbunds webbplats .
beroende på årstiden och området finns det olika aktivitetsmöjligheter .
Språkvalet kan påverka barnets möjligheter att studera olika språk i skolan .
finska som andra språk i den grundläggande undervisningenfinska _ svenska
Programguideengelska
beskattning
de inkomster som du har haft från början av året
i Finland ska man alltid på förhand komma överens om besök hos andra , även hos goda vänner .
i södra Finland reser man ibland också midsommarstången .
Socialbyråerna betjänar kommuninvånarna till exempel i följande ärenden :
medling kan ofta vara nyttig och hjälpa er att komma överens i olika frågor utan rättegång .
de har tagit lån eller finansierat sin bostad på andra sätt .
mån @-@ fre kl . 8.15 @-@ 16.00
många flygbolag erbjuder flyg från Finland till utlandet .
bevis för yrkeskunnighet med fristående examen
Väestöliittos mentorskap i fråga om arbetskarriär är avsett för utbildade invandrare .
din flytt till Finland kan betraktas som stadigvarande i följande situationer :
åldringar kan använda tjänsterna vid de vanliga hälsostationerna .
också myndigheterna måste följa lagen .
Områdeskoordinatorerfinska
möjligheter att studera finska eller svenska
när du tar hand om en gammal eller sjuk anhörig eller en anhörig med funktionsnedsättning för att han eller hon ska kunna bo kvar i sitt hem , kan du ha rätt till stöd för närståendevård .
om din bostad har skadats , till exempel till följd av brand eller vattenskada , kan hemförsäkringen i vissa fall ersätta de extra boendekostnaderna .
huruvida du behöver ett uppehållstillstånd beror på i vilket land du är medborgare , varför du kommer till Finland och hur länge du ska stanna .
be om kontaktuppgifterna till patientombudsmannen vid den vårdenhet där du har varit klient .
Skattebeloppet justeras i efterskott utgående från hur stora dina inkomster och avdrag verkligen har varit .
allmän information om studier i finska och svenska i Finland hittar du på InfoFinlands sida Finska och svenska språket .
mer information om medling i familjefrågor hittar du på InfoFinlands sida Skilsmässa .
i krigen förlorade Finland områden till Sovjetunionen .
när du är utomlands kan din sociala trygghet påverkas till exempel av att du inleder studier eller börjar arbeta .
om du är företagare kan du bli medlem i företagarnas intressebevakningsorganisation Grankulla företagare rf som erbjuder sina medlemmar utbildning , nätverk och rådgivning .
olika lån har olika villkor .
på webbtjänsten kan du söka och reservera material .
magistraten utreder om du kan få en hemkommun registrerad .
till dagvårdsplatser för verksamhetsåret som börjar i augusti ansöker man senast i slutet av mars .
handikappade barns fritid
barnet har rätt att få undervisning i sin egen religion i skolan .
Arbetspensionen intjänas med det egna lönearbetet och företagandet .
i Finland finns en lag om likabehandling , som föreskriver att arbetsgivaren ska övervaka att jämställdheten på arbetsplatsen realiseras och att ingen diskrimineras på arbetsplatsen .
tfn 045.639.6274
sexuell hälsa hos kvinnor
du kan kontakta rådgivningen via den centraliserade telefontjänsten ( 06 ) 826.4477 .
makarna kan vara partiellt vårdlediga samtidigt så att den ena förkortar sin arbetstid från morgonen och den andra från eftermiddagen .
utöver pension kan FPA betala ut bostadsbidrag till pensionstagare med låga inkomster .
på InfoFinlands sida Ansökan till utbildning finns information om hur du ansöker till utbildning på andra stadiet och högskoleutbildning i Finland .
läs mer på InfoFinlands sida Stöd för vård av barn i hemmet .
Räntestöd beviljas för unga som skaffar sin första ägarbostad .
om du har betalat för lite i skatt , blir du tvungen att betala kvarskatt ( jäännösvero ) .
förskoleundervisningen börjar i augusti och anmälan ska göras i februari .
information om kontaktuppgifter finns på Vanda stads webbplats .
i Finland är nätspänningen 230 volt .
MoniNet är ett mångkulturellt center i Rovaniemi , Lappland . det upprätthålls av föreningen Rovalan Setlementti ry .
studerande
vårdnadshavare till en finsk medborgarefinska _ svenska _ engelska
ansökan till en yrkesinriktad vuxenutbildning
information om tolktjänsterfinska
mångsidiga övningar i finska språketfinska
Grankulla stad erbjuder olika tjänster för handikappade , till exempel hjälpmedel och dagverksamhet .
läkaren skriver en remiss till det sjukhus där aborten görs .
om du behöver psykisk hjälp och psykiskt stöd kan du kontakta hälsostationen .
fysiska symptom , utan att medicinska orsaker hittas för dessa
i en del kommuner kan du delta i integrationsutbildning på svenska .
om du och din sambo är bosatta i olika stater anses gemensamt boende till exempel under semesterresor inte som en tillräcklig grund för beviljande av uppehållstillstånd .
inkomsterna för din partner som är bosatt i Finland beaktas inte .
Badhuset / + simhallen Vesihiisifinska
om du behöver rättshjälp , kan du kontakta Helsingfors rättshjälpsbyrå ( Helsingin oikeusaputoimisto ) .
medlingen är kostnadsfri .
denna gräns mellan Religionerna finns fortfarande , men med reformationen byttes den katolska tron till den lutherska .
kommunerna är skyldiga att ordna många olika tjänster för sina invånare .
var får jag hjälp ?
Vuxengymnasiumfinska
stöd och hjälp för handikappade invandrarefinska _ svenska _ engelska _ ryska _ somaliska _ persiska _ arabiska _ kurdiska
kommunerna måste tillhandahålla handikappade de tjänster som de behöver .
privata servicehusfinska
när föräldrarna har kommit överens om barnets boende , vårdnad , umgängesrätt och underhållsbidrag kan socialväsendet på orten bekräfta avtalet .
Studieutbudet är väldigt mångsidigt .
om bostaden har centralvärme , ingår uppvärmningen i allmänhet i hyran .
vid rådgivningen följs moderns , fostrets och hela familjens hälsotillstånd under graviditeten .
i anslutning till TE @-@ byrån finns ett rum där man kan uträtta ärenden på egen hand .
i Grankulla finns också privata tandläkare .
din grundutbildning avgör till hurudan yrkesutbildning du kan söka och på vilket sätt ansökan sker .
i Helsingfors , Åbo , Tammerfors och Esbo får barn och gravida kvinnor samma hälso- och sjukvårdstjänster som övriga invånare .
ekonomiskt stöd under den yrkesinriktade arbetskraftsutbildningen
till exempel finns det information om kurserna i finska språket i Helsingfors , Tammerfors och Åbo i tjänsten Finnishcourses.fi .
sexuell hälsa hos män
i Esbo finns flera bibliotek på olika håll i staden .
preventivmedel säljs på apoteket .
hur kan man minska mängden avfall ?
anmäl dig som arbetssökande i TE @-@ byråns webbtjänst .
om ett barn blir sjukt och behöver snabbt vård , ta kontakt med hälsostationen ( terveysasema ) .
många medborgarorganisationer och föreningar har särskilda ungdomsavdelningar som ordnar verksamhet för unga .
information för flyktingarfinska _ engelska _ franska _ persiska _ arabiska _ kurdiska
du kan ofta boka läkartiden via mödrarådgivningen .
självrisktiden är vanligen den dag då du insjuknade och därpå följande nio vardagar .
Finland blev självständigt 1917 .
linkkiArbets- och näringsministeriet :
följ informationen på arbetsplatsen .
om detta inte hjälper , kan du kontakta disponenten eller hyresvärden .
Serviceguide för handikappade invandrare ( pdf , 797,26 ) finska _ engelska _ ryska _ arabiska
de sköter begravningsarrangemangen , som till exempel transporten av den avlidne .
stödet är avsett för dem som har en hemkommun i Finland .
Finland har 5,5 miljoner invånare .
konflikter med grannarna
den är avsedd för de elever som ännu inte har särskilt bra kunskaper i finska .
linkkiAvfallsverksföreningen :
om du vistas utomlands tillfälligt , det vill säga under ett år , betalar FPA vanligtvis din pension som vanligt .
att studera i Finland
hyresvärden har rätt att häva hyresavtalet om du inte betalar din hyra .
att tvinga någon till äktenskap är ett brott i Finland .
Hälsostationernafinska _ svenska _ engelska
hälsostationerna har öppet från måndag till fredag , vanligen kl . 8 @-@ 16 .
kontaktuppgifter till enheten som väljer hyresgästerna , telefontid kl . 12 @-@ 15 :
om till exempel utbildning i läs- och skrivkunnighet eller någon annan språkutbildning har godkänts till din integrationsplan , tas det inte ut någon avgift för studierna .
du kan vända dig till diskrimineringsombudsmannen till exempel om du själv har råkat ut för etnisk diskriminering eller observerat att en annan person diskrimineras .
fråga din arbetsgivare som hen använder tjänsten Enter Finland för arbetsgivare .
linkkiFaro :
om din finländska arbetsgivare har sänt dig utomlands för att arbeta förlorar du inte ditt uppehållstillstånd i Finland även om du vistas utomlands på grund av arbetet i över två år .
Uleåborg
dessutom övervakar riksdagen regeringens verksamhet .
om familjen har barn under 18 år och äktenskapet slutar ska föräldrarna i samband med skilsmässan komma överens om följande :
Grankulla socialbyrå
vinterkriget och fortsättningskriget
skattebyrån , om du behöver personbeteckningen för beskattningen .
skattebyrån ( verotoimisto ) har ett serviceställe i centrala Helsingfors .
ansökan kan även göras senare , men då tillämpas kravet på tillräcklig inkomst .
vanligtvis kan man få FPA:s bidrag då de övriga inkomsterna är låga .
detta får inte orsaka extra kostnader för patienten .
när du ansöker om ditt första uppehållstillstånd i Finland kan du även be om att bli registrerad i Finlands befolkningsdatasystem .
om du har ett uppehållstillstånd för arbetstagare som endast gäller arbete för en viss arbetsgivare och du förlorar din arbetsplats , ska du ansöka om ett nytt uppehållstillstånd för arbetstagare eller ett uppehållstillstånd på andra grunder .
för att få bostadsbidrag måste du också du omfattas av den sociala tryggheten i Finland .
i vissa fall kan du alltså inte få webbankkoder även om du har ett bankkonto .
anvisningar för jobbintervjunfinska _ svenska _ engelska
du kan ansöka om finskt medborgarskap när du har fyllt 18 år , har bott permanent i Finland i tillräckligt många år , har nöjaktiga muntliga och skriftliga kunskaper i finska eller svenska eller motsvarande kunskaper i finskt eller finlandssvenskt teckenspråk och din identitet är tillförlitligt utredd .
om du inte avbokar debiteras du på en avgift om 27 euro .
barn
12 @-@ 17 år och adoptivbarn till en finsk medborgare
rehabilitering för gravt handikappade
grunderna för antagning av studeranden beror på utbildningen .
familjerådgivningfinska _ engelska
i Finland finns många patientföreningar som tillhandahåller information och rådgivning för människor med en viss sjukdom .
samtal till Nollalinja är kostnadsfria och de syns inte i telefonräkningen .
sådana stipendier är till exempel de som beviljats av staten , läroanstalter eller organisationer .
också tillräckliga medel är en grund .
föräldrapenning
Stadin aikuisopisto ordnar i vissa lekparker och familjehus kurser i finska för invandrarföräldrar .
invandrartjänster
du har ett gemensamt barn med din sambo ( då uteblir kravet på gemensamt boende under två års tid ) eller
om det finns minst tio anställda på en arbetsplats väljer dessa ut en arbetarskyddsfullmäktig som representerar dem .
vid behov skriver läkaren en remiss till den psykiatriska polikliniken för dig .
du kan även ansöka till yrkesutbildning för vuxna .
läs mer på InfoFinlands sida Gymnasieförberedande utbildning .
val av vigselform
Övernattningsalternativ i Karlebyfinska _ svenska _ engelska
modersmålsprovet är ett obligatoriskt prov i studentexamen .
privata hyresbostäder
en familjebostad är en omöblerad lägenhet som endast hyrs ut till personer i samma hushåll .
du kan grunda ett aktiebolag antingen själv eller tillsammans med andra delägare .
förmodligen får du en tid snabbare på en privat hälsostation än inom den offentliga hälsovården .
du kan också boka tid hos en privat tandläkare .
stödet kommer från samhället i form av den sociala tryggheten .
kom ihåg att kontrollera också det nya beskattningsbeslutet .
du kan utarbeta en integrationsplan t.ex. med en arbetskraftsrådgivare vid arbets- och näringsbyrån , alltså TE @-@ byrån ( TE @-@ toimisto ) , eller med en socialarbetare på socialbyrån .
du har rätt att utnyttja de offentliga hälsovårdstjänsterna om du har hemkommun i Finland .
mer information om dessa språk får du på webbplatsen för Forskningscentralen för de inhemska språken .
det är lättare att söka jobb om du vet hur en examen som du avlagt utomlands motsvarar en finländsk examen .
på InfoFinlands sida Utbildning i Grankulla finns information om dagvård för barn .
i Finland ägs cirka 70 procent av idrottsanläggningarna av kommunerna .
jag är lärare / ingenjör / studerande .
äktenskapsförord är frivilligt .
även om finländarna i allmänhet behärskar engelska relativt väl har du ändå mycket nytta av att kunna finska eller svenska .
telefon : 040.806.8101
om du inte kan betala dina räkningar eller skulder då de förfaller , ska du kontakta skuldrådgivningen ( velkaneuvonta ) .
du kan söka svenskspråkiga högskoleutbildningar via tjänsten Opintopolku.fi .
information om småbarnspedagogikfinska _ svenska _ engelska
köp endast sådana saker du behöver .
Motionsrekommendationerfinska _ engelska
om du vill förbättra dina kunskaper i finska eller svenska innan du söker till ett gymnasium , kan du söka till en förberedande gymnasieutbildning .
hjälp till diskrimineringsofferfinska _ svenska _ engelska _ ryska _ estniska _ franska _ somaliska _ spanska _ turkiska _ kinesiska _ persiska _ arabiska _ kurdiska _ albanska _ tyska _ thai _ vietnamesiska _ portugisiska _ tagalog _ polska
Studentbostäderna är oftast billigare än bostäderna på den öppna marknaden .
boka en tid på mödrarådgivningen .
Grunddagpenningfinska _ svenska _ engelska
anmäl dig till husets ägare .
en läkare eller någon annan yrkesutbildad person avgör detta .
om du behöver stöd för din integration , utarbetas en integrationsplan för dig efter den inledande kartläggningen .
observera att officiella handlingar som tagits med från utlandet ska vara legaliserade och i original samt översatta till finska , svenska eller engelska .
faderskapspenning .
privat tandvård är dyrare än offentlig tandvård .
Handikappades rättigheter
enligt Finlands lag är äktenskapet ( avioliitto ) ett lagstadgat förhållande mellan två människor .
på gymnasiet kan man även höja vitsorden i sitt avgångsbetyg eller studera enskilda ämnen .
om barnet inte kan få krävande medicinska rehabilitering från FPA , ska rehabiliteringen ordnas av hemkommunen .
att slå , sparka och knuffa
linkkiBortförda barn rf :
det självständiga Finland blev en republik där lagarna stiftas av en folkvald riksdag .
du kan även studera språket på Internet .
hälsovårdstjänster ges i Finland på finska och svenska .
om du inte har en finländsk personbeteckning , är ditt bibliotekskort i kraft ett år i taget .
Tänk på att frivilligarbete kan påverka din arbetslöshetsförsäkring .
påsen tillsluts noga .
olika läkarstationer erbjuder olika tjänster .
Förnamnen ska vara förenliga med Finlands namnlag .
information om jobbsökning i Finland hittar du på InfoFinlands sida Var hittar jag jobb ?
svenskspråkiga yrkesläroanstalter och gymnasieskolor finns i svenskspråkiga och tvåspråkiga kommuner och i en del finskspråkiga kommuner .
uppsägningstiden är den tid som arbetstagaren är skyldig att arbeta innan arbetet upphör .
boendetjänster för handikappadefinska _ svenska _ engelska
Finland ligger i Nordeuropa .
under Ryssland blev Finland ett speciellt område som utvecklades på kejsarens order .
om du vill ta en personförsäkring i ett finländskt försäkringsbolag ska du vanligtvis ha ett finländskt FPA @-@ kort .
ibland krävs att du lyckas tillräckligt bra med dina studier för att du ska få ett stipendium .
underhållsbidraget har på grund av förälderns ekonomiska situation fastställts till ett belopp som underskrider underhållsstödet .
uppehållstillstånd för studerande från andra EU @-@ länder
yrkeshögskoleexamen kan avläggas på 3,5 @-@ 4,5 år .
Helsingfors är även ett viktigt centrum för affärs- och kulturlivet .
gymnasiet ger förberedande utbildning till exempel för yrkeshögskola och universitet .
en talskada
om originalspråket för ditt betyg inte är finska , svenska eller engelska behöver du vanligtvis en officiell översättning av handlingarna som görs av en auktoriserad översättare .
vem som helst kan studera vid dessa .
information om tjänster för äldrefinska _ svenska _ engelska
det är bra att förvara filten till exempel i närheten av spisen .
inom företagshälsovården har arbetstagaren tillgång till hälsovårdarens , företagsläkarens och företagspsykologens tjänster .
om du flyttar utomlands
att låna material
om du eller din familj har utgifter på grund av särskilda behov , för vilka du inte kan få grundläggande utkomststöd , kan socialbyrån i din hemkommun bevilja kompletterande och förebyggande utkomststöd ( täydentävä ja ehkäisevä toimeentulotuki ) .
tfn 050.300.6093
om du kommer till Finland för att studera kan du få en studentbostad där du får bo så länge som dina studier i Finland pågår .
förskoleundervisningen ordnas av kommunerna och är kostnadsfri för familjen .
vård av barn
du kan rösta i kommunalvalet om :
information om diskrimineringfinska _ svenska _ engelska
Hedersrelaterat våld
att bo i en bostadsrättsbostad är ett alternativ till att köpa eller hyra sin bostad .
på beskattningen inverkar också huruvida din arbetsgivare är ett finländskt eller ett utländskt företag .
det är lättast om operationen görs innan graviditeten har börjat , men den kan också göras i mitten av graviditeten .
om du bor i östra Helsingfors , sydöstra Helsingfors , nordöstra Helsingfors eller norra Helsingfors hittar du hälsovårdscentraljouren vid Malms sjukhus .
Besläktade språk är till exempel estniska och ungerska .
Besöksadress :
Fennovoima bygger kärnkraftverksenheten Hanhikivi 1 i Pyhäjoki .
Helsingfors stad hjälper arbetslösa helsingforsare att hitta jobb eller utbildning .
vid social delaktighet ,
du kan byta ut ditt körkort till ett finskt körkort på Ajovarmas serviceställe .
barnet kan också få hjälpmedel om han eller hon inte kan studera utan dem eller om det är mycket svårt utan dem .
att bevittna våldsamma situationer
om du redan har fött fyra barn
stödet består antingen av pengar eller tjänster .
Vinter
lönen kan innehålla olika förmåner .
du är medborgare i ett nordiskt land
om du misstänker att du har en könssjukdom kan du boka en läkartid på hälsostationen eller en privat läkarstation .
Finskans uttal är mycket regelbundet .
sådana är till exempel många idrotts- och simhallar och andra idrottsanläggningar , såsom fotbollsplaner och skridskobanor .
du kan själv välja om du vill ta ut 25 procent eller 50 procent av beloppet på din månatliga arbetspension .
om du behöver mer information om legalisering av handlingar , kontakta magistraten eller utrikesministeriet i ditt eget land .
för att få en inledande kartläggning gjord , ska du anmäla dig som arbetssökande via Internet på adressen te @-@ palvelut.fi .
prepaid @-@ kortet är i förväg laddat med en summa som man sedan kan ringa för .
dessa uppgifter är bland annat namn , födelsedatum , medborgarskap , kön och adress .
fler än 400.000 finländare lämnade de förlorade områdena och kom som flyktingar till övriga delar av landet .
i Kelviå , ca 10 km norrut från Karleby , finns Toivonen djurpark och drängmuseum .
anmäl diskrimineringfinska _ svenska _ engelska
verksamheten i öppna daghem och invånarparker är kostnadsfri och du behöver inte anmäla dig på förhand .
du kan ändå behöva ett visum .
läs mera om privatvårdsstöd på Fpa:s sidor .
andra religiösa samfund i Finland är till exempel katolska kyrkan i Finland , Pingstkyrkan i Finland , Frikyrkan i Finland , Adventkyrkan i Finland , mormonkyrkan och Jehovas vittnen .
IHH - serviceställe för dig som flyttar till Finland engelska
du ska vanligtvis även kunna visa ditt betalningsbeteende , dvs. uppgifter som visar att du har betalat dina räkningar och inte har några betalningsanmärkningar .
det är tillåtet att spela in material på offentliga platser , för inspelning i privata lokaler ska tillstånd inhämtas .
föreningens styrelse
Borgmästaren och stadens aktörer ordnar boendemöten runtom i Helsingfors för invånarna där man berättar om och diskuterar stadens ärenden .
vem som helst kan studera vid en öppen högskola .
Förvara hyresavtalet noga .
öppna linjen : 09.7562.2260
hjälp för unga
